//32x32 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 922 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize,base_dat_a,base_dat_b,cpu_addr; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [4:0]regaddr1,regaddr2,rdata,adata; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
wire hht;
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 

control t1 (Clk,base_dat_a,base_dat_b,addr1,addr2,dataIn1,dataIn2,Rst,RD,csize,cpu_addr,hht,regaddr1,regaddr2,rdata,adata);


initial begin 
Clk = 1'b0; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1;
cpu_addr = 32'd126;
  v_values_base = 32'd2; 
  matrix_base = 32'd170 ; 
  wdata_col_base = 32'd10920 ; 
  row_base = 32'd118420 ; 
  csize = COL_SIZE; 
  //fe_init = 1'b0; 
// RD = 1'b0; 
// RD = 1'b1; 
 #99600; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 

if(regaddr1 == 5'd6)
	base_dat_a = wdata_col_base;
else if (regaddr1 == 5'd8)
	base_dat_a = v_values_base;

if(regaddr2 == 5'd15) begin
	base_dat_b = row_base; 
 end
else if (regaddr2 == 5'd9)
	base_dat_b = matrix_base;

case(addr1)  
32'd118420: dataIn1 = 32'd0
; 
32'd118421: dataIn1 = 32'd26
; 
32'd118422: dataIn1 = 32'd51
; 
32'd118423: dataIn1 = 32'd80
; 
32'd118424: dataIn1 = 32'd107
; 
32'd118425: dataIn1 = 32'd133
; 
32'd118426: dataIn1 = 32'd161
; 
32'd118427: dataIn1 = 32'd187
; 
32'd118428: dataIn1 = 32'd214
; 
32'd118429: dataIn1 = 32'd242
; 
32'd118430: dataIn1 = 32'd270
; 
32'd118431: dataIn1 = 32'd297
; 
32'd118432: dataIn1 = 32'd326
; 
32'd118433: dataIn1 = 32'd354
; 
32'd118434: dataIn1 = 32'd379
; 
32'd118435: dataIn1 = 32'd409
; 
32'd118436: dataIn1 = 32'd436
; 
32'd118437: dataIn1 = 32'd463
; 
32'd118438: dataIn1 = 32'd489
; 
32'd118439: dataIn1 = 32'd515
; 
32'd118440: dataIn1 = 32'd539
; 
32'd118441: dataIn1 = 32'd568
; 
32'd118442: dataIn1 = 32'd595
; 
32'd118443: dataIn1 = 32'd624
; 
32'd118444: dataIn1 = 32'd653
; 
32'd118445: dataIn1 = 32'd679
; 
32'd118446: dataIn1 = 32'd708
; 
32'd118447: dataIn1 = 32'd733
; 
32'd118448: dataIn1 = 32'd763
; 
32'd118449: dataIn1 = 32'd789
; 
32'd118450: dataIn1 = 32'd816
; 
32'd118451: dataIn1 = 32'd842
; 
32'd118452: dataIn1 = 32'd868
; 
32'd10920: dataIn1 = 32'd0
; 
32'd10921: dataIn1 = 32'd26
; 
32'd10922: dataIn1 = 32'd51
; 
32'd10923: dataIn1 = 32'd80
; 
32'd10924: dataIn1 = 32'd107
; 
32'd10925: dataIn1 = 32'd133
; 
32'd10926: dataIn1 = 32'd161
; 
32'd10927: dataIn1 = 32'd187
; 
32'd10928: dataIn1 = 32'd214
; 
32'd10929: dataIn1 = 32'd242
; 
32'd10930: dataIn1 = 32'd270
; 
32'd10931: dataIn1 = 32'd297
; 
32'd10932: dataIn1 = 32'd326
; 
32'd10933: dataIn1 = 32'd354
; 
32'd10934: dataIn1 = 32'd379
; 
32'd10935: dataIn1 = 32'd409
; 
32'd10936: dataIn1 = 32'd436
; 
32'd10937: dataIn1 = 32'd463
; 
32'd10938: dataIn1 = 32'd489
; 
32'd10939: dataIn1 = 32'd515
; 
32'd10940: dataIn1 = 32'd539
; 
32'd10941: dataIn1 = 32'd568
; 
32'd10942: dataIn1 = 32'd595
; 
32'd10943: dataIn1 = 32'd624
; 
32'd10944: dataIn1 = 32'd653
; 
32'd10945: dataIn1 = 32'd679
; 
32'd10946: dataIn1 = 32'd708
; 
32'd10947: dataIn1 = 32'd733
; 
32'd10948: dataIn1 = 32'd763
; 
32'd10949: dataIn1 = 32'd789
; 
32'd10950: dataIn1 = 32'd816
; 
32'd10951: dataIn1 = 32'd842
; 
32'd10952: dataIn1 = 32'd868
; 
32'd10953: dataIn1 = 32'd1
; 
32'd10954: dataIn1 = 32'd3
; 
32'd10955: dataIn1 = 32'd4
; 
32'd10956: dataIn1 = 32'd5
; 
32'd10957: dataIn1 = 32'd6
; 
32'd10958: dataIn1 = 32'd8
; 
32'd10959: dataIn1 = 32'd9
; 
32'd10960: dataIn1 = 32'd10
; 
32'd10961: dataIn1 = 32'd11
; 
32'd10962: dataIn1 = 32'd12
; 
32'd10963: dataIn1 = 32'd13
; 
32'd10964: dataIn1 = 32'd14
; 
32'd10965: dataIn1 = 32'd15
; 
32'd10966: dataIn1 = 32'd16
; 
32'd10967: dataIn1 = 32'd17
; 
32'd10968: dataIn1 = 32'd18
; 
32'd10969: dataIn1 = 32'd20
; 
32'd10970: dataIn1 = 32'd22
; 
32'd10971: dataIn1 = 32'd23
; 
32'd10972: dataIn1 = 32'd24
; 
32'd10973: dataIn1 = 32'd25
; 
32'd10974: dataIn1 = 32'd26
; 
32'd10975: dataIn1 = 32'd27
; 
32'd10976: dataIn1 = 32'd28
; 
32'd10977: dataIn1 = 32'd29
; 
32'd10978: dataIn1 = 32'd31
; 
32'd10979: dataIn1 = 32'd0
; 
32'd10980: dataIn1 = 32'd1
; 
32'd10981: dataIn1 = 32'd2
; 
32'd10982: dataIn1 = 32'd3
; 
32'd10983: dataIn1 = 32'd4
; 
32'd10984: dataIn1 = 32'd6
; 
32'd10985: dataIn1 = 32'd8
; 
32'd10986: dataIn1 = 32'd9
; 
32'd10987: dataIn1 = 32'd11
; 
32'd10988: dataIn1 = 32'd12
; 
32'd10989: dataIn1 = 32'd13
; 
32'd10990: dataIn1 = 32'd15
; 
32'd10991: dataIn1 = 32'd16
; 
32'd10992: dataIn1 = 32'd17
; 
32'd10993: dataIn1 = 32'd20
; 
32'd10994: dataIn1 = 32'd21
; 
32'd10995: dataIn1 = 32'd22
; 
32'd10996: dataIn1 = 32'd23
; 
32'd10997: dataIn1 = 32'd24
; 
32'd10998: dataIn1 = 32'd25
; 
32'd10999: dataIn1 = 32'd26
; 
32'd11000: dataIn1 = 32'd28
; 
32'd11001: dataIn1 = 32'd29
; 
32'd11002: dataIn1 = 32'd30
; 
32'd11003: dataIn1 = 32'd31
; 
32'd11004: dataIn1 = 32'd0
; 
32'd11005: dataIn1 = 32'd1
; 
32'd11006: dataIn1 = 32'd2
; 
32'd11007: dataIn1 = 32'd3
; 
32'd11008: dataIn1 = 32'd4
; 
32'd11009: dataIn1 = 32'd5
; 
32'd11010: dataIn1 = 32'd6
; 
32'd11011: dataIn1 = 32'd7
; 
32'd11012: dataIn1 = 32'd8
; 
32'd11013: dataIn1 = 32'd9
; 
32'd11014: dataIn1 = 32'd10
; 
32'd11015: dataIn1 = 32'd11
; 
32'd11016: dataIn1 = 32'd12
; 
32'd11017: dataIn1 = 32'd13
; 
32'd11018: dataIn1 = 32'd14
; 
32'd11019: dataIn1 = 32'd16
; 
32'd11020: dataIn1 = 32'd17
; 
32'd11021: dataIn1 = 32'd18
; 
32'd11022: dataIn1 = 32'd20
; 
32'd11023: dataIn1 = 32'd21
; 
32'd11024: dataIn1 = 32'd23
; 
32'd11025: dataIn1 = 32'd24
; 
32'd11026: dataIn1 = 32'd25
; 
32'd11027: dataIn1 = 32'd26
; 
32'd11028: dataIn1 = 32'd27
; 
32'd11029: dataIn1 = 32'd28
; 
32'd11030: dataIn1 = 32'd29
; 
32'd11031: dataIn1 = 32'd30
; 
32'd11032: dataIn1 = 32'd31
; 
32'd11033: dataIn1 = 32'd0
; 
32'd11034: dataIn1 = 32'd1
; 
32'd11035: dataIn1 = 32'd2
; 
32'd11036: dataIn1 = 32'd3
; 
32'd11037: dataIn1 = 32'd5
; 
32'd11038: dataIn1 = 32'd6
; 
32'd11039: dataIn1 = 32'd7
; 
32'd11040: dataIn1 = 32'd8
; 
32'd11041: dataIn1 = 32'd10
; 
32'd11042: dataIn1 = 32'd12
; 
32'd11043: dataIn1 = 32'd13
; 
32'd11044: dataIn1 = 32'd14
; 
32'd11045: dataIn1 = 32'd15
; 
32'd11046: dataIn1 = 32'd16
; 
32'd11047: dataIn1 = 32'd17
; 
32'd11048: dataIn1 = 32'd18
; 
32'd11049: dataIn1 = 32'd19
; 
32'd11050: dataIn1 = 32'd20
; 
32'd11051: dataIn1 = 32'd21
; 
32'd11052: dataIn1 = 32'd22
; 
32'd11053: dataIn1 = 32'd25
; 
32'd11054: dataIn1 = 32'd26
; 
32'd11055: dataIn1 = 32'd27
; 
32'd11056: dataIn1 = 32'd28
; 
32'd11057: dataIn1 = 32'd29
; 
32'd11058: dataIn1 = 32'd30
; 
32'd11059: dataIn1 = 32'd31
; 
32'd11060: dataIn1 = 32'd1
; 
32'd11061: dataIn1 = 32'd2
; 
32'd11062: dataIn1 = 32'd4
; 
32'd11063: dataIn1 = 32'd5
; 
32'd11064: dataIn1 = 32'd6
; 
32'd11065: dataIn1 = 32'd7
; 
32'd11066: dataIn1 = 32'd8
; 
32'd11067: dataIn1 = 32'd10
; 
32'd11068: dataIn1 = 32'd11
; 
32'd11069: dataIn1 = 32'd12
; 
32'd11070: dataIn1 = 32'd14
; 
32'd11071: dataIn1 = 32'd15
; 
32'd11072: dataIn1 = 32'd16
; 
32'd11073: dataIn1 = 32'd17
; 
32'd11074: dataIn1 = 32'd18
; 
32'd11075: dataIn1 = 32'd19
; 
32'd11076: dataIn1 = 32'd20
; 
32'd11077: dataIn1 = 32'd21
; 
32'd11078: dataIn1 = 32'd22
; 
32'd11079: dataIn1 = 32'd23
; 
32'd11080: dataIn1 = 32'd24
; 
32'd11081: dataIn1 = 32'd26
; 
32'd11082: dataIn1 = 32'd27
; 
32'd11083: dataIn1 = 32'd28
; 
32'd11084: dataIn1 = 32'd29
; 
32'd11085: dataIn1 = 32'd30
; 
32'd11086: dataIn1 = 32'd0
; 
32'd11087: dataIn1 = 32'd2
; 
32'd11088: dataIn1 = 32'd3
; 
32'd11089: dataIn1 = 32'd4
; 
32'd11090: dataIn1 = 32'd5
; 
32'd11091: dataIn1 = 32'd6
; 
32'd11092: dataIn1 = 32'd7
; 
32'd11093: dataIn1 = 32'd8
; 
32'd11094: dataIn1 = 32'd10
; 
32'd11095: dataIn1 = 32'd11
; 
32'd11096: dataIn1 = 32'd12
; 
32'd11097: dataIn1 = 32'd13
; 
32'd11098: dataIn1 = 32'd14
; 
32'd11099: dataIn1 = 32'd15
; 
32'd11100: dataIn1 = 32'd17
; 
32'd11101: dataIn1 = 32'd18
; 
32'd11102: dataIn1 = 32'd19
; 
32'd11103: dataIn1 = 32'd20
; 
32'd11104: dataIn1 = 32'd21
; 
32'd11105: dataIn1 = 32'd22
; 
32'd11106: dataIn1 = 32'd23
; 
32'd11107: dataIn1 = 32'd24
; 
32'd11108: dataIn1 = 32'd25
; 
32'd11109: dataIn1 = 32'd26
; 
32'd11110: dataIn1 = 32'd28
; 
32'd11111: dataIn1 = 32'd29
; 
32'd11112: dataIn1 = 32'd30
; 
32'd11113: dataIn1 = 32'd31
; 
32'd11114: dataIn1 = 32'd0
; 
32'd11115: dataIn1 = 32'd1
; 
32'd11116: dataIn1 = 32'd2
; 
32'd11117: dataIn1 = 32'd3
; 
32'd11118: dataIn1 = 32'd4
; 
32'd11119: dataIn1 = 32'd6
; 
32'd11120: dataIn1 = 32'd7
; 
32'd11121: dataIn1 = 32'd9
; 
32'd11122: dataIn1 = 32'd10
; 
32'd11123: dataIn1 = 32'd11
; 
32'd11124: dataIn1 = 32'd12
; 
32'd11125: dataIn1 = 32'd13
; 
32'd11126: dataIn1 = 32'd14
; 
32'd11127: dataIn1 = 32'd15
; 
32'd11128: dataIn1 = 32'd16
; 
32'd11129: dataIn1 = 32'd18
; 
32'd11130: dataIn1 = 32'd20
; 
32'd11131: dataIn1 = 32'd22
; 
32'd11132: dataIn1 = 32'd23
; 
32'd11133: dataIn1 = 32'd24
; 
32'd11134: dataIn1 = 32'd25
; 
32'd11135: dataIn1 = 32'd26
; 
32'd11136: dataIn1 = 32'd28
; 
32'd11137: dataIn1 = 32'd29
; 
32'd11138: dataIn1 = 32'd30
; 
32'd11139: dataIn1 = 32'd31
; 
32'd11140: dataIn1 = 32'd0
; 
32'd11141: dataIn1 = 32'd1
; 
32'd11142: dataIn1 = 32'd2
; 
32'd11143: dataIn1 = 32'd3
; 
32'd11144: dataIn1 = 32'd4
; 
32'd11145: dataIn1 = 32'd5
; 
32'd11146: dataIn1 = 32'd6
; 
32'd11147: dataIn1 = 32'd7
; 
32'd11148: dataIn1 = 32'd8
; 
32'd11149: dataIn1 = 32'd9
; 
32'd11150: dataIn1 = 32'd11
; 
32'd11151: dataIn1 = 32'd12
; 
32'd11152: dataIn1 = 32'd13
; 
32'd11153: dataIn1 = 32'd14
; 
32'd11154: dataIn1 = 32'd15
; 
32'd11155: dataIn1 = 32'd16
; 
32'd11156: dataIn1 = 32'd17
; 
32'd11157: dataIn1 = 32'd18
; 
32'd11158: dataIn1 = 32'd21
; 
32'd11159: dataIn1 = 32'd22
; 
32'd11160: dataIn1 = 32'd23
; 
32'd11161: dataIn1 = 32'd24
; 
32'd11162: dataIn1 = 32'd26
; 
32'd11163: dataIn1 = 32'd27
; 
32'd11164: dataIn1 = 32'd29
; 
32'd11165: dataIn1 = 32'd30
; 
32'd11166: dataIn1 = 32'd31
; 
32'd11167: dataIn1 = 32'd1
; 
32'd11168: dataIn1 = 32'd2
; 
32'd11169: dataIn1 = 32'd3
; 
32'd11170: dataIn1 = 32'd4
; 
32'd11171: dataIn1 = 32'd5
; 
32'd11172: dataIn1 = 32'd6
; 
32'd11173: dataIn1 = 32'd7
; 
32'd11174: dataIn1 = 32'd8
; 
32'd11175: dataIn1 = 32'd9
; 
32'd11176: dataIn1 = 32'd10
; 
32'd11177: dataIn1 = 32'd11
; 
32'd11178: dataIn1 = 32'd12
; 
32'd11179: dataIn1 = 32'd13
; 
32'd11180: dataIn1 = 32'd14
; 
32'd11181: dataIn1 = 32'd15
; 
32'd11182: dataIn1 = 32'd16
; 
32'd11183: dataIn1 = 32'd17
; 
32'd11184: dataIn1 = 32'd18
; 
32'd11185: dataIn1 = 32'd19
; 
32'd11186: dataIn1 = 32'd21
; 
32'd11187: dataIn1 = 32'd22
; 
32'd11188: dataIn1 = 32'd23
; 
32'd11189: dataIn1 = 32'd26
; 
32'd11190: dataIn1 = 32'd27
; 
32'd11191: dataIn1 = 32'd28
; 
32'd11192: dataIn1 = 32'd29
; 
32'd11193: dataIn1 = 32'd30
; 
32'd11194: dataIn1 = 32'd31
; 
32'd11195: dataIn1 = 32'd0
; 
32'd11196: dataIn1 = 32'd1
; 
32'd11197: dataIn1 = 32'd2
; 
32'd11198: dataIn1 = 32'd3
; 
32'd11199: dataIn1 = 32'd4
; 
32'd11200: dataIn1 = 32'd5
; 
32'd11201: dataIn1 = 32'd6
; 
32'd11202: dataIn1 = 32'd7
; 
32'd11203: dataIn1 = 32'd9
; 
32'd11204: dataIn1 = 32'd10
; 
32'd11205: dataIn1 = 32'd11
; 
32'd11206: dataIn1 = 32'd12
; 
32'd11207: dataIn1 = 32'd13
; 
32'd11208: dataIn1 = 32'd14
; 
32'd11209: dataIn1 = 32'd15
; 
32'd11210: dataIn1 = 32'd17
; 
32'd11211: dataIn1 = 32'd18
; 
32'd11212: dataIn1 = 32'd20
; 
32'd11213: dataIn1 = 32'd21
; 
32'd11214: dataIn1 = 32'd22
; 
32'd11215: dataIn1 = 32'd23
; 
32'd11216: dataIn1 = 32'd24
; 
32'd11217: dataIn1 = 32'd25
; 
32'd11218: dataIn1 = 32'd26
; 
32'd11219: dataIn1 = 32'd27
; 
32'd11220: dataIn1 = 32'd28
; 
32'd11221: dataIn1 = 32'd29
; 
32'd11222: dataIn1 = 32'd30
; 
32'd11223: dataIn1 = 32'd0
; 
32'd11224: dataIn1 = 32'd1
; 
32'd11225: dataIn1 = 32'd2
; 
32'd11226: dataIn1 = 32'd3
; 
32'd11227: dataIn1 = 32'd4
; 
32'd11228: dataIn1 = 32'd5
; 
32'd11229: dataIn1 = 32'd6
; 
32'd11230: dataIn1 = 32'd7
; 
32'd11231: dataIn1 = 32'd8
; 
32'd11232: dataIn1 = 32'd9
; 
32'd11233: dataIn1 = 32'd10
; 
32'd11234: dataIn1 = 32'd11
; 
32'd11235: dataIn1 = 32'd13
; 
32'd11236: dataIn1 = 32'd14
; 
32'd11237: dataIn1 = 32'd15
; 
32'd11238: dataIn1 = 32'd16
; 
32'd11239: dataIn1 = 32'd18
; 
32'd11240: dataIn1 = 32'd19
; 
32'd11241: dataIn1 = 32'd20
; 
32'd11242: dataIn1 = 32'd23
; 
32'd11243: dataIn1 = 32'd24
; 
32'd11244: dataIn1 = 32'd25
; 
32'd11245: dataIn1 = 32'd26
; 
32'd11246: dataIn1 = 32'd27
; 
32'd11247: dataIn1 = 32'd28
; 
32'd11248: dataIn1 = 32'd29
; 
32'd11249: dataIn1 = 32'd31
; 
32'd11250: dataIn1 = 32'd0
; 
32'd11251: dataIn1 = 32'd1
; 
32'd11252: dataIn1 = 32'd2
; 
32'd11253: dataIn1 = 32'd3
; 
32'd11254: dataIn1 = 32'd4
; 
32'd11255: dataIn1 = 32'd5
; 
32'd11256: dataIn1 = 32'd6
; 
32'd11257: dataIn1 = 32'd7
; 
32'd11258: dataIn1 = 32'd8
; 
32'd11259: dataIn1 = 32'd9
; 
32'd11260: dataIn1 = 32'd10
; 
32'd11261: dataIn1 = 32'd11
; 
32'd11262: dataIn1 = 32'd12
; 
32'd11263: dataIn1 = 32'd13
; 
32'd11264: dataIn1 = 32'd14
; 
32'd11265: dataIn1 = 32'd15
; 
32'd11266: dataIn1 = 32'd16
; 
32'd11267: dataIn1 = 32'd17
; 
32'd11268: dataIn1 = 32'd18
; 
32'd11269: dataIn1 = 32'd19
; 
32'd11270: dataIn1 = 32'd22
; 
32'd11271: dataIn1 = 32'd23
; 
32'd11272: dataIn1 = 32'd24
; 
32'd11273: dataIn1 = 32'd25
; 
32'd11274: dataIn1 = 32'd26
; 
32'd11275: dataIn1 = 32'd27
; 
32'd11276: dataIn1 = 32'd28
; 
32'd11277: dataIn1 = 32'd29
; 
32'd11278: dataIn1 = 32'd31
; 
32'd11279: dataIn1 = 32'd0
; 
32'd11280: dataIn1 = 32'd2
; 
32'd11281: dataIn1 = 32'd3
; 
32'd11282: dataIn1 = 32'd4
; 
32'd11283: dataIn1 = 32'd5
; 
32'd11284: dataIn1 = 32'd6
; 
32'd11285: dataIn1 = 32'd7
; 
32'd11286: dataIn1 = 32'd8
; 
32'd11287: dataIn1 = 32'd9
; 
32'd11288: dataIn1 = 32'd10
; 
32'd11289: dataIn1 = 32'd11
; 
32'd11290: dataIn1 = 32'd12
; 
32'd11291: dataIn1 = 32'd13
; 
32'd11292: dataIn1 = 32'd14
; 
32'd11293: dataIn1 = 32'd16
; 
32'd11294: dataIn1 = 32'd17
; 
32'd11295: dataIn1 = 32'd18
; 
32'd11296: dataIn1 = 32'd19
; 
32'd11297: dataIn1 = 32'd20
; 
32'd11298: dataIn1 = 32'd22
; 
32'd11299: dataIn1 = 32'd23
; 
32'd11300: dataIn1 = 32'd24
; 
32'd11301: dataIn1 = 32'd25
; 
32'd11302: dataIn1 = 32'd26
; 
32'd11303: dataIn1 = 32'd27
; 
32'd11304: dataIn1 = 32'd28
; 
32'd11305: dataIn1 = 32'd30
; 
32'd11306: dataIn1 = 32'd31
; 
32'd11307: dataIn1 = 32'd0
; 
32'd11308: dataIn1 = 32'd1
; 
32'd11309: dataIn1 = 32'd2
; 
32'd11310: dataIn1 = 32'd4
; 
32'd11311: dataIn1 = 32'd5
; 
32'd11312: dataIn1 = 32'd7
; 
32'd11313: dataIn1 = 32'd8
; 
32'd11314: dataIn1 = 32'd9
; 
32'd11315: dataIn1 = 32'd10
; 
32'd11316: dataIn1 = 32'd11
; 
32'd11317: dataIn1 = 32'd12
; 
32'd11318: dataIn1 = 32'd13
; 
32'd11319: dataIn1 = 32'd14
; 
32'd11320: dataIn1 = 32'd15
; 
32'd11321: dataIn1 = 32'd17
; 
32'd11322: dataIn1 = 32'd18
; 
32'd11323: dataIn1 = 32'd19
; 
32'd11324: dataIn1 = 32'd20
; 
32'd11325: dataIn1 = 32'd22
; 
32'd11326: dataIn1 = 32'd23
; 
32'd11327: dataIn1 = 32'd25
; 
32'd11328: dataIn1 = 32'd26
; 
32'd11329: dataIn1 = 32'd27
; 
32'd11330: dataIn1 = 32'd28
; 
32'd11331: dataIn1 = 32'd30
; 
32'd11332: dataIn1 = 32'd0
; 
32'd11333: dataIn1 = 32'd1
; 
32'd11334: dataIn1 = 32'd2
; 
32'd11335: dataIn1 = 32'd3
; 
32'd11336: dataIn1 = 32'd4
; 
32'd11337: dataIn1 = 32'd5
; 
32'd11338: dataIn1 = 32'd6
; 
32'd11339: dataIn1 = 32'd7
; 
32'd11340: dataIn1 = 32'd8
; 
32'd11341: dataIn1 = 32'd9
; 
32'd11342: dataIn1 = 32'd10
; 
32'd11343: dataIn1 = 32'd11
; 
32'd11344: dataIn1 = 32'd12
; 
32'd11345: dataIn1 = 32'd14
; 
32'd11346: dataIn1 = 32'd16
; 
32'd11347: dataIn1 = 32'd17
; 
32'd11348: dataIn1 = 32'd18
; 
32'd11349: dataIn1 = 32'd19
; 
32'd11350: dataIn1 = 32'd20
; 
32'd11351: dataIn1 = 32'd21
; 
32'd11352: dataIn1 = 32'd22
; 
32'd11353: dataIn1 = 32'd23
; 
32'd11354: dataIn1 = 32'd24
; 
32'd11355: dataIn1 = 32'd25
; 
32'd11356: dataIn1 = 32'd26
; 
32'd11357: dataIn1 = 32'd27
; 
32'd11358: dataIn1 = 32'd28
; 
32'd11359: dataIn1 = 32'd29
; 
32'd11360: dataIn1 = 32'd30
; 
32'd11361: dataIn1 = 32'd31
; 
32'd11362: dataIn1 = 32'd0
; 
32'd11363: dataIn1 = 32'd1
; 
32'd11364: dataIn1 = 32'd2
; 
32'd11365: dataIn1 = 32'd3
; 
32'd11366: dataIn1 = 32'd5
; 
32'd11367: dataIn1 = 32'd6
; 
32'd11368: dataIn1 = 32'd7
; 
32'd11369: dataIn1 = 32'd8
; 
32'd11370: dataIn1 = 32'd9
; 
32'd11371: dataIn1 = 32'd10
; 
32'd11372: dataIn1 = 32'd11
; 
32'd11373: dataIn1 = 32'd12
; 
32'd11374: dataIn1 = 32'd13
; 
32'd11375: dataIn1 = 32'd14
; 
32'd11376: dataIn1 = 32'd15
; 
32'd11377: dataIn1 = 32'd17
; 
32'd11378: dataIn1 = 32'd18
; 
32'd11379: dataIn1 = 32'd20
; 
32'd11380: dataIn1 = 32'd21
; 
32'd11381: dataIn1 = 32'd23
; 
32'd11382: dataIn1 = 32'd24
; 
32'd11383: dataIn1 = 32'd25
; 
32'd11384: dataIn1 = 32'd26
; 
32'd11385: dataIn1 = 32'd27
; 
32'd11386: dataIn1 = 32'd28
; 
32'd11387: dataIn1 = 32'd29
; 
32'd11388: dataIn1 = 32'd30
; 
32'd11389: dataIn1 = 32'd0
; 
32'd11390: dataIn1 = 32'd1
; 
32'd11391: dataIn1 = 32'd2
; 
32'd11392: dataIn1 = 32'd4
; 
32'd11393: dataIn1 = 32'd5
; 
32'd11394: dataIn1 = 32'd6
; 
32'd11395: dataIn1 = 32'd7
; 
32'd11396: dataIn1 = 32'd8
; 
32'd11397: dataIn1 = 32'd9
; 
32'd11398: dataIn1 = 32'd10
; 
32'd11399: dataIn1 = 32'd11
; 
32'd11400: dataIn1 = 32'd12
; 
32'd11401: dataIn1 = 32'd13
; 
32'd11402: dataIn1 = 32'd14
; 
32'd11403: dataIn1 = 32'd15
; 
32'd11404: dataIn1 = 32'd17
; 
32'd11405: dataIn1 = 32'd18
; 
32'd11406: dataIn1 = 32'd20
; 
32'd11407: dataIn1 = 32'd21
; 
32'd11408: dataIn1 = 32'd22
; 
32'd11409: dataIn1 = 32'd23
; 
32'd11410: dataIn1 = 32'd25
; 
32'd11411: dataIn1 = 32'd26
; 
32'd11412: dataIn1 = 32'd27
; 
32'd11413: dataIn1 = 32'd28
; 
32'd11414: dataIn1 = 32'd30
; 
32'd11415: dataIn1 = 32'd31
; 
32'd11416: dataIn1 = 32'd0
; 
32'd11417: dataIn1 = 32'd1
; 
32'd11418: dataIn1 = 32'd2
; 
32'd11419: dataIn1 = 32'd3
; 
32'd11420: dataIn1 = 32'd4
; 
32'd11421: dataIn1 = 32'd5
; 
32'd11422: dataIn1 = 32'd6
; 
32'd11423: dataIn1 = 32'd7
; 
32'd11424: dataIn1 = 32'd8
; 
32'd11425: dataIn1 = 32'd9
; 
32'd11426: dataIn1 = 32'd10
; 
32'd11427: dataIn1 = 32'd11
; 
32'd11428: dataIn1 = 32'd12
; 
32'd11429: dataIn1 = 32'd13
; 
32'd11430: dataIn1 = 32'd14
; 
32'd11431: dataIn1 = 32'd16
; 
32'd11432: dataIn1 = 32'd17
; 
32'd11433: dataIn1 = 32'd18
; 
32'd11434: dataIn1 = 32'd20
; 
32'd11435: dataIn1 = 32'd22
; 
32'd11436: dataIn1 = 32'd24
; 
32'd11437: dataIn1 = 32'd25
; 
32'd11438: dataIn1 = 32'd26
; 
32'd11439: dataIn1 = 32'd28
; 
32'd11440: dataIn1 = 32'd29
; 
32'd11441: dataIn1 = 32'd31
; 
32'd11442: dataIn1 = 32'd0
; 
32'd11443: dataIn1 = 32'd1
; 
32'd11444: dataIn1 = 32'd2
; 
32'd11445: dataIn1 = 32'd3
; 
32'd11446: dataIn1 = 32'd4
; 
32'd11447: dataIn1 = 32'd5
; 
32'd11448: dataIn1 = 32'd6
; 
32'd11449: dataIn1 = 32'd8
; 
32'd11450: dataIn1 = 32'd9
; 
32'd11451: dataIn1 = 32'd10
; 
32'd11452: dataIn1 = 32'd12
; 
32'd11453: dataIn1 = 32'd13
; 
32'd11454: dataIn1 = 32'd14
; 
32'd11455: dataIn1 = 32'd15
; 
32'd11456: dataIn1 = 32'd17
; 
32'd11457: dataIn1 = 32'd18
; 
32'd11458: dataIn1 = 32'd19
; 
32'd11459: dataIn1 = 32'd20
; 
32'd11460: dataIn1 = 32'd23
; 
32'd11461: dataIn1 = 32'd24
; 
32'd11462: dataIn1 = 32'd25
; 
32'd11463: dataIn1 = 32'd26
; 
32'd11464: dataIn1 = 32'd27
; 
32'd11465: dataIn1 = 32'd29
; 
32'd11466: dataIn1 = 32'd30
; 
32'd11467: dataIn1 = 32'd31
; 
32'd11468: dataIn1 = 32'd0
; 
32'd11469: dataIn1 = 32'd2
; 
32'd11470: dataIn1 = 32'd4
; 
32'd11471: dataIn1 = 32'd5
; 
32'd11472: dataIn1 = 32'd7
; 
32'd11473: dataIn1 = 32'd8
; 
32'd11474: dataIn1 = 32'd10
; 
32'd11475: dataIn1 = 32'd11
; 
32'd11476: dataIn1 = 32'd12
; 
32'd11477: dataIn1 = 32'd13
; 
32'd11478: dataIn1 = 32'd14
; 
32'd11479: dataIn1 = 32'd15
; 
32'd11480: dataIn1 = 32'd16
; 
32'd11481: dataIn1 = 32'd18
; 
32'd11482: dataIn1 = 32'd21
; 
32'd11483: dataIn1 = 32'd22
; 
32'd11484: dataIn1 = 32'd23
; 
32'd11485: dataIn1 = 32'd24
; 
32'd11486: dataIn1 = 32'd25
; 
32'd11487: dataIn1 = 32'd26
; 
32'd11488: dataIn1 = 32'd27
; 
32'd11489: dataIn1 = 32'd28
; 
32'd11490: dataIn1 = 32'd29
; 
32'd11491: dataIn1 = 32'd30
; 
32'd11492: dataIn1 = 32'd0
; 
32'd11493: dataIn1 = 32'd1
; 
32'd11494: dataIn1 = 32'd2
; 
32'd11495: dataIn1 = 32'd4
; 
32'd11496: dataIn1 = 32'd5
; 
32'd11497: dataIn1 = 32'd6
; 
32'd11498: dataIn1 = 32'd8
; 
32'd11499: dataIn1 = 32'd9
; 
32'd11500: dataIn1 = 32'd10
; 
32'd11501: dataIn1 = 32'd11
; 
32'd11502: dataIn1 = 32'd12
; 
32'd11503: dataIn1 = 32'd13
; 
32'd11504: dataIn1 = 32'd14
; 
32'd11505: dataIn1 = 32'd16
; 
32'd11506: dataIn1 = 32'd17
; 
32'd11507: dataIn1 = 32'd18
; 
32'd11508: dataIn1 = 32'd19
; 
32'd11509: dataIn1 = 32'd20
; 
32'd11510: dataIn1 = 32'd21
; 
32'd11511: dataIn1 = 32'd22
; 
32'd11512: dataIn1 = 32'd23
; 
32'd11513: dataIn1 = 32'd24
; 
32'd11514: dataIn1 = 32'd25
; 
32'd11515: dataIn1 = 32'd26
; 
32'd11516: dataIn1 = 32'd27
; 
32'd11517: dataIn1 = 32'd28
; 
32'd11518: dataIn1 = 32'd29
; 
32'd11519: dataIn1 = 32'd30
; 
32'd11520: dataIn1 = 32'd31
; 
32'd11521: dataIn1 = 32'd1
; 
32'd11522: dataIn1 = 32'd2
; 
32'd11523: dataIn1 = 32'd3
; 
32'd11524: dataIn1 = 32'd4
; 
32'd11525: dataIn1 = 32'd6
; 
32'd11526: dataIn1 = 32'd7
; 
32'd11527: dataIn1 = 32'd8
; 
32'd11528: dataIn1 = 32'd9
; 
32'd11529: dataIn1 = 32'd10
; 
32'd11530: dataIn1 = 32'd11
; 
32'd11531: dataIn1 = 32'd12
; 
32'd11532: dataIn1 = 32'd13
; 
32'd11533: dataIn1 = 32'd14
; 
32'd11534: dataIn1 = 32'd15
; 
32'd11535: dataIn1 = 32'd16
; 
32'd11536: dataIn1 = 32'd17
; 
32'd11537: dataIn1 = 32'd18
; 
32'd11538: dataIn1 = 32'd20
; 
32'd11539: dataIn1 = 32'd21
; 
32'd11540: dataIn1 = 32'd22
; 
32'd11541: dataIn1 = 32'd24
; 
32'd11542: dataIn1 = 32'd26
; 
32'd11543: dataIn1 = 32'd27
; 
32'd11544: dataIn1 = 32'd28
; 
32'd11545: dataIn1 = 32'd29
; 
32'd11546: dataIn1 = 32'd30
; 
32'd11547: dataIn1 = 32'd31
; 
32'd11548: dataIn1 = 32'd0
; 
32'd11549: dataIn1 = 32'd1
; 
32'd11550: dataIn1 = 32'd2
; 
32'd11551: dataIn1 = 32'd3
; 
32'd11552: dataIn1 = 32'd4
; 
32'd11553: dataIn1 = 32'd5
; 
32'd11554: dataIn1 = 32'd6
; 
32'd11555: dataIn1 = 32'd7
; 
32'd11556: dataIn1 = 32'd8
; 
32'd11557: dataIn1 = 32'd9
; 
32'd11558: dataIn1 = 32'd10
; 
32'd11559: dataIn1 = 32'd11
; 
32'd11560: dataIn1 = 32'd12
; 
32'd11561: dataIn1 = 32'd14
; 
32'd11562: dataIn1 = 32'd15
; 
32'd11563: dataIn1 = 32'd16
; 
32'd11564: dataIn1 = 32'd18
; 
32'd11565: dataIn1 = 32'd19
; 
32'd11566: dataIn1 = 32'd20
; 
32'd11567: dataIn1 = 32'd21
; 
32'd11568: dataIn1 = 32'd23
; 
32'd11569: dataIn1 = 32'd24
; 
32'd11570: dataIn1 = 32'd25
; 
32'd11571: dataIn1 = 32'd26
; 
32'd11572: dataIn1 = 32'd27
; 
32'd11573: dataIn1 = 32'd28
; 
32'd11574: dataIn1 = 32'd29
; 
32'd11575: dataIn1 = 32'd30
; 
32'd11576: dataIn1 = 32'd31
; 
32'd11577: dataIn1 = 32'd1
; 
32'd11578: dataIn1 = 32'd2
; 
32'd11579: dataIn1 = 32'd3
; 
32'd11580: dataIn1 = 32'd4
; 
32'd11581: dataIn1 = 32'd5
; 
32'd11582: dataIn1 = 32'd6
; 
32'd11583: dataIn1 = 32'd7
; 
32'd11584: dataIn1 = 32'd8
; 
32'd11585: dataIn1 = 32'd9
; 
32'd11586: dataIn1 = 32'd11
; 
32'd11587: dataIn1 = 32'd12
; 
32'd11588: dataIn1 = 32'd13
; 
32'd11589: dataIn1 = 32'd14
; 
32'd11590: dataIn1 = 32'd15
; 
32'd11591: dataIn1 = 32'd16
; 
32'd11592: dataIn1 = 32'd17
; 
32'd11593: dataIn1 = 32'd18
; 
32'd11594: dataIn1 = 32'd19
; 
32'd11595: dataIn1 = 32'd20
; 
32'd11596: dataIn1 = 32'd21
; 
32'd11597: dataIn1 = 32'd23
; 
32'd11598: dataIn1 = 32'd24
; 
32'd11599: dataIn1 = 32'd25
; 
32'd11600: dataIn1 = 32'd26
; 
32'd11601: dataIn1 = 32'd27
; 
32'd11602: dataIn1 = 32'd28
; 
32'd11603: dataIn1 = 32'd29
; 
32'd11604: dataIn1 = 32'd30
; 
32'd11605: dataIn1 = 32'd31
; 
32'd11606: dataIn1 = 32'd0
; 
32'd11607: dataIn1 = 32'd1
; 
32'd11608: dataIn1 = 32'd2
; 
32'd11609: dataIn1 = 32'd3
; 
32'd11610: dataIn1 = 32'd6
; 
32'd11611: dataIn1 = 32'd7
; 
32'd11612: dataIn1 = 32'd8
; 
32'd11613: dataIn1 = 32'd9
; 
32'd11614: dataIn1 = 32'd10
; 
32'd11615: dataIn1 = 32'd11
; 
32'd11616: dataIn1 = 32'd12
; 
32'd11617: dataIn1 = 32'd13
; 
32'd11618: dataIn1 = 32'd14
; 
32'd11619: dataIn1 = 32'd16
; 
32'd11620: dataIn1 = 32'd17
; 
32'd11621: dataIn1 = 32'd18
; 
32'd11622: dataIn1 = 32'd19
; 
32'd11623: dataIn1 = 32'd20
; 
32'd11624: dataIn1 = 32'd21
; 
32'd11625: dataIn1 = 32'd22
; 
32'd11626: dataIn1 = 32'd23
; 
32'd11627: dataIn1 = 32'd24
; 
32'd11628: dataIn1 = 32'd25
; 
32'd11629: dataIn1 = 32'd27
; 
32'd11630: dataIn1 = 32'd28
; 
32'd11631: dataIn1 = 32'd29
; 
32'd11632: dataIn1 = 32'd0
; 
32'd11633: dataIn1 = 32'd1
; 
32'd11634: dataIn1 = 32'd2
; 
32'd11635: dataIn1 = 32'd3
; 
32'd11636: dataIn1 = 32'd4
; 
32'd11637: dataIn1 = 32'd5
; 
32'd11638: dataIn1 = 32'd6
; 
32'd11639: dataIn1 = 32'd7
; 
32'd11640: dataIn1 = 32'd8
; 
32'd11641: dataIn1 = 32'd9
; 
32'd11642: dataIn1 = 32'd10
; 
32'd11643: dataIn1 = 32'd11
; 
32'd11644: dataIn1 = 32'd12
; 
32'd11645: dataIn1 = 32'd13
; 
32'd11646: dataIn1 = 32'd14
; 
32'd11647: dataIn1 = 32'd15
; 
32'd11648: dataIn1 = 32'd16
; 
32'd11649: dataIn1 = 32'd17
; 
32'd11650: dataIn1 = 32'd19
; 
32'd11651: dataIn1 = 32'd20
; 
32'd11652: dataIn1 = 32'd21
; 
32'd11653: dataIn1 = 32'd22
; 
32'd11654: dataIn1 = 32'd24
; 
32'd11655: dataIn1 = 32'd25
; 
32'd11656: dataIn1 = 32'd26
; 
32'd11657: dataIn1 = 32'd27
; 
32'd11658: dataIn1 = 32'd28
; 
32'd11659: dataIn1 = 32'd29
; 
32'd11660: dataIn1 = 32'd30
; 
32'd11661: dataIn1 = 32'd0
; 
32'd11662: dataIn1 = 32'd1
; 
32'd11663: dataIn1 = 32'd4
; 
32'd11664: dataIn1 = 32'd5
; 
32'd11665: dataIn1 = 32'd6
; 
32'd11666: dataIn1 = 32'd7
; 
32'd11667: dataIn1 = 32'd9
; 
32'd11668: dataIn1 = 32'd12
; 
32'd11669: dataIn1 = 32'd13
; 
32'd11670: dataIn1 = 32'd14
; 
32'd11671: dataIn1 = 32'd15
; 
32'd11672: dataIn1 = 32'd16
; 
32'd11673: dataIn1 = 32'd17
; 
32'd11674: dataIn1 = 32'd18
; 
32'd11675: dataIn1 = 32'd19
; 
32'd11676: dataIn1 = 32'd21
; 
32'd11677: dataIn1 = 32'd22
; 
32'd11678: dataIn1 = 32'd23
; 
32'd11679: dataIn1 = 32'd24
; 
32'd11680: dataIn1 = 32'd26
; 
32'd11681: dataIn1 = 32'd27
; 
32'd11682: dataIn1 = 32'd28
; 
32'd11683: dataIn1 = 32'd29
; 
32'd11684: dataIn1 = 32'd30
; 
32'd11685: dataIn1 = 32'd31
; 
32'd11686: dataIn1 = 32'd0
; 
32'd11687: dataIn1 = 32'd1
; 
32'd11688: dataIn1 = 32'd2
; 
32'd11689: dataIn1 = 32'd3
; 
32'd11690: dataIn1 = 32'd4
; 
32'd11691: dataIn1 = 32'd5
; 
32'd11692: dataIn1 = 32'd7
; 
32'd11693: dataIn1 = 32'd8
; 
32'd11694: dataIn1 = 32'd9
; 
32'd11695: dataIn1 = 32'd10
; 
32'd11696: dataIn1 = 32'd11
; 
32'd11697: dataIn1 = 32'd12
; 
32'd11698: dataIn1 = 32'd13
; 
32'd11699: dataIn1 = 32'd14
; 
32'd11700: dataIn1 = 32'd15
; 
32'd11701: dataIn1 = 32'd16
; 
32'd11702: dataIn1 = 32'd17
; 
32'd11703: dataIn1 = 32'd18
; 
32'd11704: dataIn1 = 32'd19
; 
32'd11705: dataIn1 = 32'd20
; 
32'd11706: dataIn1 = 32'd21
; 
32'd11707: dataIn1 = 32'd22
; 
32'd11708: dataIn1 = 32'd23
; 
32'd11709: dataIn1 = 32'd24
; 
32'd11710: dataIn1 = 32'd25
; 
32'd11711: dataIn1 = 32'd27
; 
32'd11712: dataIn1 = 32'd28
; 
32'd11713: dataIn1 = 32'd29
; 
32'd11714: dataIn1 = 32'd30
; 
32'd11715: dataIn1 = 32'd31
; 
32'd11716: dataIn1 = 32'd0
; 
32'd11717: dataIn1 = 32'd1
; 
32'd11718: dataIn1 = 32'd2
; 
32'd11719: dataIn1 = 32'd3
; 
32'd11720: dataIn1 = 32'd4
; 
32'd11721: dataIn1 = 32'd5
; 
32'd11722: dataIn1 = 32'd6
; 
32'd11723: dataIn1 = 32'd7
; 
32'd11724: dataIn1 = 32'd8
; 
32'd11725: dataIn1 = 32'd9
; 
32'd11726: dataIn1 = 32'd12
; 
32'd11727: dataIn1 = 32'd14
; 
32'd11728: dataIn1 = 32'd15
; 
32'd11729: dataIn1 = 32'd16
; 
32'd11730: dataIn1 = 32'd17
; 
32'd11731: dataIn1 = 32'd18
; 
32'd11732: dataIn1 = 32'd19
; 
32'd11733: dataIn1 = 32'd21
; 
32'd11734: dataIn1 = 32'd22
; 
32'd11735: dataIn1 = 32'd23
; 
32'd11736: dataIn1 = 32'd24
; 
32'd11737: dataIn1 = 32'd25
; 
32'd11738: dataIn1 = 32'd26
; 
32'd11739: dataIn1 = 32'd27
; 
32'd11740: dataIn1 = 32'd29
; 
32'd11741: dataIn1 = 32'd30
; 
32'd11742: dataIn1 = 32'd0
; 
32'd11743: dataIn1 = 32'd1
; 
32'd11744: dataIn1 = 32'd2
; 
32'd11745: dataIn1 = 32'd3
; 
32'd11746: dataIn1 = 32'd4
; 
32'd11747: dataIn1 = 32'd6
; 
32'd11748: dataIn1 = 32'd7
; 
32'd11749: dataIn1 = 32'd8
; 
32'd11750: dataIn1 = 32'd9
; 
32'd11751: dataIn1 = 32'd10
; 
32'd11752: dataIn1 = 32'd11
; 
32'd11753: dataIn1 = 32'd12
; 
32'd11754: dataIn1 = 32'd14
; 
32'd11755: dataIn1 = 32'd15
; 
32'd11756: dataIn1 = 32'd16
; 
32'd11757: dataIn1 = 32'd17
; 
32'd11758: dataIn1 = 32'd18
; 
32'd11759: dataIn1 = 32'd20
; 
32'd11760: dataIn1 = 32'd21
; 
32'd11761: dataIn1 = 32'd22
; 
32'd11762: dataIn1 = 32'd23
; 
32'd11763: dataIn1 = 32'd26
; 
32'd11764: dataIn1 = 32'd27
; 
32'd11765: dataIn1 = 32'd28
; 
32'd11766: dataIn1 = 32'd29
; 
32'd11767: dataIn1 = 32'd30
; 
32'd11768: dataIn1 = 32'd31
; 
32'd11769: dataIn1 = 32'd0
; 
32'd11770: dataIn1 = 32'd1
; 
32'd11771: dataIn1 = 32'd2
; 
32'd11772: dataIn1 = 32'd3
; 
32'd11773: dataIn1 = 32'd4
; 
32'd11774: dataIn1 = 32'd5
; 
32'd11775: dataIn1 = 32'd6
; 
32'd11776: dataIn1 = 32'd7
; 
32'd11777: dataIn1 = 32'd8
; 
32'd11778: dataIn1 = 32'd9
; 
32'd11779: dataIn1 = 32'd10
; 
32'd11780: dataIn1 = 32'd12
; 
32'd11781: dataIn1 = 32'd13
; 
32'd11782: dataIn1 = 32'd15
; 
32'd11783: dataIn1 = 32'd17
; 
32'd11784: dataIn1 = 32'd18
; 
32'd11785: dataIn1 = 32'd19
; 
32'd11786: dataIn1 = 32'd20
; 
32'd11787: dataIn1 = 32'd22
; 
32'd11788: dataIn1 = 32'd23
; 
32'd11789: dataIn1 = 32'd24
; 
32'd11790: dataIn1 = 32'd25
; 
32'd11791: dataIn1 = 32'd26
; 
32'd11792: dataIn1 = 32'd27
; 
32'd11793: dataIn1 = 32'd29
; 
32'd11794: dataIn1 = 32'd30
; 
32'd11795: dataIn1 = 32'd0
; 
32'd11796: dataIn1 = 32'd1
; 
32'd11797: dataIn1 = 32'd2
; 
32'd11798: dataIn1 = 32'd3
; 
32'd11799: dataIn1 = 32'd4
; 
32'd11800: dataIn1 = 32'd5
; 
32'd11801: dataIn1 = 32'd6
; 
32'd11802: dataIn1 = 32'd7
; 
32'd11803: dataIn1 = 32'd8
; 
32'd11804: dataIn1 = 32'd9
; 
32'd11805: dataIn1 = 32'd11
; 
32'd11806: dataIn1 = 32'd12
; 
32'd11807: dataIn1 = 32'd14
; 
32'd11808: dataIn1 = 32'd18
; 
32'd11809: dataIn1 = 32'd19
; 
32'd11810: dataIn1 = 32'd20
; 
32'd11811: dataIn1 = 32'd21
; 
32'd11812: dataIn1 = 32'd23
; 
32'd11813: dataIn1 = 32'd24
; 
32'd11814: dataIn1 = 32'd25
; 
32'd11815: dataIn1 = 32'd26
; 
32'd11816: dataIn1 = 32'd27
; 
32'd11817: dataIn1 = 32'd28
; 
32'd11818: dataIn1 = 32'd29
; 
32'd11819: dataIn1 = 32'd30
; 
32'd11820: dataIn1 = 32'd31
; 
32'd11821: dataIn1 = 32'd0; 
32'd11822: dataIn1 = 32'd1; 
32'd11823: dataIn1 = 32'd2; 
32'd11824: dataIn1 = 32'd3; 
32'd11825: dataIn1 = 32'd4; 
32'd11826: dataIn1 = 32'd5; 
32'd11827: dataIn1 = 32'd6; 
32'd11828: dataIn1 = 32'd7; 
32'd11829: dataIn1 = 32'd8; 
32'd11830: dataIn1 = 32'd9; 
32'd11831: dataIn1 = 32'd10; 
32'd11832: dataIn1 = 32'd11; 
32'd11833: dataIn1 = 32'd12; 
32'd11834: dataIn1 = 32'd13; 
32'd11835: dataIn1 = 32'd14; 
32'd11836: dataIn1 = 32'd15; 
32'd11837: dataIn1 = 32'd16; 
32'd11838: dataIn1 = 32'd17; 
32'd11839: dataIn1 = 32'd18; 
32'd11840: dataIn1 = 32'd19; 
32'd11841: dataIn1 = 32'd20; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd11; 
32'd3: dataIn2 = 32'd98; 
32'd4: dataIn2 = 32'd45; 
32'd5: dataIn2 = 32'd53; 
32'd6: dataIn2 = 32'd75; 
32'd7: dataIn2 = 32'd67; 
32'd8: dataIn2 = 32'd26; 
32'd9: dataIn2 = 32'd40; 
32'd10: dataIn2 = 32'd47; 
32'd11: dataIn2 = 32'd35; 
32'd12: dataIn2 = 32'd39; 
32'd13: dataIn2 = 32'd51; 
32'd14: dataIn2 = 32'd57; 
32'd15: dataIn2 = 32'd11; 
32'd16: dataIn2 = 32'd51; 
32'd17: dataIn2 = 32'd74; 
32'd18: dataIn2 = 32'd65; 
32'd19: dataIn2 = 32'd56; 
32'd20: dataIn2 = 32'd90; 
32'd21: dataIn2 = 32'd43; 
32'd22: dataIn2 = 32'd85; 
32'd23: dataIn2 = 32'd19; 
32'd24: dataIn2 = 32'd68; 
32'd25: dataIn2 = 32'd14; 
32'd26: dataIn2 = 32'd82; 
32'd27: dataIn2 = 32'd79; 
32'd28: dataIn2 = 32'd12; 
32'd29: dataIn2 = 32'd1; 
32'd30: dataIn2 = 32'd15; 
32'd31: dataIn2 = 32'd27; 
32'd32: dataIn2 = 32'd77; 
32'd33: dataIn2 = 32'd51; 
default: 
	dataIn2 = 32'd99999; 
endcase 
case(addr2) 

32'd170: dataIn2 = 32'd50; 
32'd171: dataIn2 = 32'd3; 
32'd172: dataIn2 = 32'd94; 
32'd173: dataIn2 = 32'd34; 
32'd174: dataIn2 = 32'd23; 
32'd175: dataIn2 = 32'd89; 
32'd176: dataIn2 = 32'd6; 
32'd177: dataIn2 = 32'd80; 
32'd178: dataIn2 = 32'd90; 
32'd179: dataIn2 = 32'd34; 
32'd180: dataIn2 = 32'd46; 
32'd181: dataIn2 = 32'd69; 
32'd182: dataIn2 = 32'd68; 
32'd183: dataIn2 = 32'd82; 
32'd184: dataIn2 = 32'd13; 
32'd185: dataIn2 = 32'd58; 
32'd186: dataIn2 = 32'd60; 
32'd187: dataIn2 = 32'd63; 
32'd188: dataIn2 = 32'd93; 
32'd189: dataIn2 = 32'd86; 
32'd190: dataIn2 = 32'd92; 
32'd191: dataIn2 = 32'd78; 
32'd192: dataIn2 = 32'd48; 
32'd193: dataIn2 = 32'd78; 
32'd194: dataIn2 = 32'd80; 
32'd195: dataIn2 = 32'd10; 
32'd196: dataIn2 = 32'd49; 
32'd197: dataIn2 = 32'd89; 
32'd198: dataIn2 = 32'd34; 
32'd199: dataIn2 = 32'd13; 
32'd200: dataIn2 = 32'd86; 
32'd201: dataIn2 = 32'd4; 
32'd202: dataIn2 = 32'd77; 
32'd203: dataIn2 = 32'd12; 
32'd204: dataIn2 = 32'd47; 
32'd205: dataIn2 = 32'd36; 
32'd206: dataIn2 = 32'd29; 
32'd207: dataIn2 = 32'd49; 
32'd208: dataIn2 = 32'd30; 
32'd209: dataIn2 = 32'd12; 
32'd210: dataIn2 = 32'd20; 
32'd211: dataIn2 = 32'd19; 
32'd212: dataIn2 = 32'd93; 
32'd213: dataIn2 = 32'd75; 
32'd214: dataIn2 = 32'd66; 
32'd215: dataIn2 = 32'd91; 
32'd216: dataIn2 = 32'd23; 
32'd217: dataIn2 = 32'd95; 
32'd218: dataIn2 = 32'd98; 
32'd219: dataIn2 = 32'd23; 
32'd220: dataIn2 = 32'd58; 
32'd221: dataIn2 = 32'd37; 
32'd222: dataIn2 = 32'd6; 
32'd223: dataIn2 = 32'd72; 
32'd224: dataIn2 = 32'd45; 
32'd225: dataIn2 = 32'd17; 
32'd226: dataIn2 = 32'd44; 
32'd227: dataIn2 = 32'd24; 
32'd228: dataIn2 = 32'd59; 
32'd229: dataIn2 = 32'd62; 
32'd230: dataIn2 = 32'd3; 
32'd231: dataIn2 = 32'd30; 
32'd232: dataIn2 = 32'd47; 
32'd233: dataIn2 = 32'd61; 
32'd234: dataIn2 = 32'd16; 
32'd235: dataIn2 = 32'd40; 
32'd236: dataIn2 = 32'd55; 
32'd237: dataIn2 = 32'd60; 
32'd238: dataIn2 = 32'd2; 
32'd239: dataIn2 = 32'd21; 
32'd240: dataIn2 = 32'd17; 
32'd241: dataIn2 = 32'd7; 
32'd242: dataIn2 = 32'd83; 
32'd243: dataIn2 = 32'd91; 
32'd244: dataIn2 = 32'd68; 
32'd245: dataIn2 = 32'd29; 
32'd246: dataIn2 = 32'd7; 
32'd247: dataIn2 = 32'd95; 
32'd248: dataIn2 = 32'd82; 
32'd249: dataIn2 = 32'd95; 
32'd250: dataIn2 = 32'd84; 
32'd251: dataIn2 = 32'd48; 
32'd252: dataIn2 = 32'd68; 
32'd253: dataIn2 = 32'd63; 
32'd254: dataIn2 = 32'd98; 
32'd255: dataIn2 = 32'd22; 
32'd256: dataIn2 = 32'd38; 
32'd257: dataIn2 = 32'd81; 
32'd258: dataIn2 = 32'd0; 
32'd259: dataIn2 = 32'd17; 
32'd260: dataIn2 = 32'd35; 
32'd261: dataIn2 = 32'd59; 
32'd262: dataIn2 = 32'd83; 
32'd263: dataIn2 = 32'd73; 
32'd264: dataIn2 = 32'd66; 
32'd265: dataIn2 = 32'd26; 
32'd266: dataIn2 = 32'd3; 
32'd267: dataIn2 = 32'd57; 
32'd268: dataIn2 = 32'd94; 
32'd269: dataIn2 = 32'd10; 
32'd270: dataIn2 = 32'd52; 
32'd271: dataIn2 = 32'd66; 
32'd272: dataIn2 = 32'd44; 
32'd273: dataIn2 = 32'd85; 
32'd274: dataIn2 = 32'd53; 
32'd275: dataIn2 = 32'd99; 
32'd276: dataIn2 = 32'd68; 
32'd277: dataIn2 = 32'd10; 
32'd278: dataIn2 = 32'd3; 
32'd279: dataIn2 = 32'd29; 
32'd280: dataIn2 = 32'd53; 
32'd281: dataIn2 = 32'd90; 
32'd282: dataIn2 = 32'd9; 
32'd283: dataIn2 = 32'd88; 
32'd284: dataIn2 = 32'd61; 
32'd285: dataIn2 = 32'd83; 
32'd286: dataIn2 = 32'd34; 
32'd287: dataIn2 = 32'd13; 
32'd288: dataIn2 = 32'd43; 
32'd289: dataIn2 = 32'd53; 
32'd290: dataIn2 = 32'd75; 
32'd291: dataIn2 = 32'd62; 
32'd292: dataIn2 = 32'd65; 
32'd293: dataIn2 = 32'd39; 
32'd294: dataIn2 = 32'd29; 
32'd295: dataIn2 = 32'd15; 
32'd296: dataIn2 = 32'd1; 
32'd297: dataIn2 = 32'd63; 
32'd298: dataIn2 = 32'd21; 
32'd299: dataIn2 = 32'd19; 
32'd300: dataIn2 = 32'd98; 
32'd301: dataIn2 = 32'd81; 
32'd302: dataIn2 = 32'd75; 
32'd303: dataIn2 = 32'd76; 
32'd304: dataIn2 = 32'd73; 
32'd305: dataIn2 = 32'd15; 
32'd306: dataIn2 = 32'd46; 
32'd307: dataIn2 = 32'd97; 
32'd308: dataIn2 = 32'd31; 
32'd309: dataIn2 = 32'd12; 
32'd310: dataIn2 = 32'd36; 
32'd311: dataIn2 = 32'd90; 
32'd312: dataIn2 = 32'd64; 
32'd313: dataIn2 = 32'd21; 
32'd314: dataIn2 = 32'd10; 
32'd315: dataIn2 = 32'd86; 
32'd316: dataIn2 = 32'd0; 
32'd317: dataIn2 = 32'd57; 
32'd318: dataIn2 = 32'd24; 
32'd319: dataIn2 = 32'd27; 
32'd320: dataIn2 = 32'd0; 
32'd321: dataIn2 = 32'd13; 
32'd322: dataIn2 = 32'd46; 
32'd323: dataIn2 = 32'd98; 
32'd324: dataIn2 = 32'd42; 
32'd325: dataIn2 = 32'd2; 
32'd326: dataIn2 = 32'd36; 
32'd327: dataIn2 = 32'd22; 
32'd328: dataIn2 = 32'd65; 
32'd329: dataIn2 = 32'd7; 
32'd330: dataIn2 = 32'd61; 
32'd331: dataIn2 = 32'd55; 
32'd332: dataIn2 = 32'd88; 
32'd333: dataIn2 = 32'd5; 
32'd334: dataIn2 = 32'd80; 
32'd335: dataIn2 = 32'd19; 
32'd336: dataIn2 = 32'd28; 
32'd337: dataIn2 = 32'd98; 
32'd338: dataIn2 = 32'd35; 
32'd339: dataIn2 = 32'd26; 
32'd340: dataIn2 = 32'd64; 
32'd341: dataIn2 = 32'd59; 
32'd342: dataIn2 = 32'd0; 
32'd343: dataIn2 = 32'd76; 
32'd344: dataIn2 = 32'd26; 
32'd345: dataIn2 = 32'd98; 
32'd346: dataIn2 = 32'd42; 
32'd347: dataIn2 = 32'd97; 
32'd348: dataIn2 = 32'd36; 
32'd349: dataIn2 = 32'd32; 
32'd350: dataIn2 = 32'd100; 
32'd351: dataIn2 = 32'd43; 
32'd352: dataIn2 = 32'd38; 
32'd353: dataIn2 = 32'd97; 
32'd354: dataIn2 = 32'd21; 
32'd355: dataIn2 = 32'd96; 
32'd356: dataIn2 = 32'd7; 
32'd357: dataIn2 = 32'd97; 
32'd358: dataIn2 = 32'd77; 
32'd359: dataIn2 = 32'd44; 
32'd360: dataIn2 = 32'd93; 
32'd361: dataIn2 = 32'd4; 
32'd362: dataIn2 = 32'd90; 
32'd363: dataIn2 = 32'd21; 
32'd364: dataIn2 = 32'd76; 
32'd365: dataIn2 = 32'd59; 
32'd366: dataIn2 = 32'd73; 
32'd367: dataIn2 = 32'd67; 
32'd368: dataIn2 = 32'd77; 
32'd369: dataIn2 = 32'd39; 
32'd370: dataIn2 = 32'd18; 
32'd371: dataIn2 = 32'd74; 
32'd372: dataIn2 = 32'd66; 
32'd373: dataIn2 = 32'd67; 
32'd374: dataIn2 = 32'd90; 
32'd375: dataIn2 = 32'd70; 
32'd376: dataIn2 = 32'd9; 
32'd377: dataIn2 = 32'd12; 
32'd378: dataIn2 = 32'd43; 
32'd379: dataIn2 = 32'd17; 
32'd380: dataIn2 = 32'd72; 
32'd381: dataIn2 = 32'd76; 
32'd382: dataIn2 = 32'd81; 
32'd383: dataIn2 = 32'd89; 
32'd384: dataIn2 = 32'd19; 
32'd385: dataIn2 = 32'd67; 
32'd386: dataIn2 = 32'd19; 
32'd387: dataIn2 = 32'd38; 
32'd388: dataIn2 = 32'd76; 
32'd389: dataIn2 = 32'd84; 
32'd390: dataIn2 = 32'd84; 
32'd391: dataIn2 = 32'd1; 
32'd392: dataIn2 = 32'd68; 
32'd393: dataIn2 = 32'd24; 
32'd394: dataIn2 = 32'd34; 
32'd395: dataIn2 = 32'd3; 
32'd396: dataIn2 = 32'd33; 
32'd397: dataIn2 = 32'd48; 
32'd398: dataIn2 = 32'd20; 
32'd399: dataIn2 = 32'd36; 
32'd400: dataIn2 = 32'd23; 
32'd401: dataIn2 = 32'd76; 
32'd402: dataIn2 = 32'd17; 
32'd403: dataIn2 = 32'd29; 
32'd404: dataIn2 = 32'd72; 
32'd405: dataIn2 = 32'd18; 
32'd406: dataIn2 = 32'd4; 
32'd407: dataIn2 = 32'd99; 
32'd408: dataIn2 = 32'd36; 
32'd409: dataIn2 = 32'd44; 
32'd410: dataIn2 = 32'd71; 
32'd411: dataIn2 = 32'd22; 
32'd412: dataIn2 = 32'd0; 
32'd413: dataIn2 = 32'd67; 
32'd414: dataIn2 = 32'd57; 
32'd415: dataIn2 = 32'd24; 
32'd416: dataIn2 = 32'd90; 
32'd417: dataIn2 = 32'd94; 
32'd418: dataIn2 = 32'd85; 
32'd419: dataIn2 = 32'd69; 
32'd420: dataIn2 = 32'd21; 
32'd421: dataIn2 = 32'd64; 
32'd422: dataIn2 = 32'd22; 
32'd423: dataIn2 = 32'd95; 
32'd424: dataIn2 = 32'd0; 
32'd425: dataIn2 = 32'd6; 
32'd426: dataIn2 = 32'd27; 
32'd427: dataIn2 = 32'd39; 
32'd428: dataIn2 = 32'd22; 
32'd429: dataIn2 = 32'd46; 
32'd430: dataIn2 = 32'd58; 
32'd431: dataIn2 = 32'd64; 
32'd432: dataIn2 = 32'd67; 
32'd433: dataIn2 = 32'd64; 
32'd434: dataIn2 = 32'd33; 
32'd435: dataIn2 = 32'd95; 
32'd436: dataIn2 = 32'd10; 
32'd437: dataIn2 = 32'd3; 
32'd438: dataIn2 = 32'd70; 
32'd439: dataIn2 = 32'd31; 
32'd440: dataIn2 = 32'd55; 
32'd441: dataIn2 = 32'd62; 
32'd442: dataIn2 = 32'd80; 
32'd443: dataIn2 = 32'd0; 
32'd444: dataIn2 = 32'd65; 
32'd445: dataIn2 = 32'd96; 
32'd446: dataIn2 = 32'd52; 
32'd447: dataIn2 = 32'd15; 
32'd448: dataIn2 = 32'd30; 
32'd449: dataIn2 = 32'd91; 
32'd450: dataIn2 = 32'd48; 
32'd451: dataIn2 = 32'd79; 
32'd452: dataIn2 = 32'd87; 
32'd453: dataIn2 = 32'd69; 
32'd454: dataIn2 = 32'd25; 
32'd455: dataIn2 = 32'd46; 
32'd456: dataIn2 = 32'd70; 
32'd457: dataIn2 = 32'd31; 
32'd458: dataIn2 = 32'd62; 
32'd459: dataIn2 = 32'd90; 
32'd460: dataIn2 = 32'd56; 
32'd461: dataIn2 = 32'd56; 
32'd462: dataIn2 = 32'd5; 
32'd463: dataIn2 = 32'd1; 
32'd464: dataIn2 = 32'd69; 
32'd465: dataIn2 = 32'd90; 
32'd466: dataIn2 = 32'd68; 
32'd467: dataIn2 = 32'd6; 
32'd468: dataIn2 = 32'd10; 
32'd469: dataIn2 = 32'd73; 
32'd470: dataIn2 = 32'd63; 
32'd471: dataIn2 = 32'd49; 
32'd472: dataIn2 = 32'd50; 
32'd473: dataIn2 = 32'd28; 
32'd474: dataIn2 = 32'd37; 
32'd475: dataIn2 = 32'd38; 
32'd476: dataIn2 = 32'd57; 
32'd477: dataIn2 = 32'd24; 
32'd478: dataIn2 = 32'd73; 
32'd479: dataIn2 = 32'd92; 
32'd480: dataIn2 = 32'd34; 
32'd481: dataIn2 = 32'd13; 
32'd482: dataIn2 = 32'd96; 
32'd483: dataIn2 = 32'd4; 
32'd484: dataIn2 = 32'd55; 
32'd485: dataIn2 = 32'd96; 
32'd486: dataIn2 = 32'd20; 
32'd487: dataIn2 = 32'd77; 
32'd488: dataIn2 = 32'd59; 
32'd489: dataIn2 = 32'd83; 
32'd490: dataIn2 = 32'd18; 
32'd491: dataIn2 = 32'd63; 
32'd492: dataIn2 = 32'd0; 
32'd493: dataIn2 = 32'd69; 
32'd494: dataIn2 = 32'd70; 
32'd495: dataIn2 = 32'd10; 
32'd496: dataIn2 = 32'd98; 
32'd497: dataIn2 = 32'd96; 
32'd498: dataIn2 = 32'd86; 
32'd499: dataIn2 = 32'd30; 
32'd500: dataIn2 = 32'd27; 
32'd501: dataIn2 = 32'd34; 
32'd502: dataIn2 = 32'd5; 
32'd503: dataIn2 = 32'd35; 
32'd504: dataIn2 = 32'd55; 
32'd505: dataIn2 = 32'd8; 
32'd506: dataIn2 = 32'd90; 
32'd507: dataIn2 = 32'd59; 
32'd508: dataIn2 = 32'd39; 
32'd509: dataIn2 = 32'd77; 
32'd510: dataIn2 = 32'd26; 
32'd511: dataIn2 = 32'd44; 
32'd512: dataIn2 = 32'd52; 
32'd513: dataIn2 = 32'd25; 
32'd514: dataIn2 = 32'd9; 
32'd515: dataIn2 = 32'd27; 
32'd516: dataIn2 = 32'd26; 
32'd517: dataIn2 = 32'd72; 
32'd518: dataIn2 = 32'd18; 
32'd519: dataIn2 = 32'd34; 
32'd520: dataIn2 = 32'd81; 
32'd521: dataIn2 = 32'd86; 
32'd522: dataIn2 = 32'd59; 
32'd523: dataIn2 = 32'd8; 
32'd524: dataIn2 = 32'd1; 
32'd525: dataIn2 = 32'd40; 
32'd526: dataIn2 = 32'd51; 
32'd527: dataIn2 = 32'd14; 
32'd528: dataIn2 = 32'd29; 
32'd529: dataIn2 = 32'd66; 
32'd530: dataIn2 = 32'd9; 
32'd531: dataIn2 = 32'd62; 
32'd532: dataIn2 = 32'd88; 
32'd533: dataIn2 = 32'd77; 
32'd534: dataIn2 = 32'd19; 
32'd535: dataIn2 = 32'd93; 
32'd536: dataIn2 = 32'd48; 
32'd537: dataIn2 = 32'd12; 
32'd538: dataIn2 = 32'd43; 
32'd539: dataIn2 = 32'd98; 
32'd540: dataIn2 = 32'd65; 
32'd541: dataIn2 = 32'd26; 
32'd542: dataIn2 = 32'd41; 
32'd543: dataIn2 = 32'd14; 
32'd544: dataIn2 = 32'd90; 
32'd545: dataIn2 = 32'd14; 
32'd546: dataIn2 = 32'd12; 
32'd547: dataIn2 = 32'd62; 
32'd548: dataIn2 = 32'd58; 
32'd549: dataIn2 = 32'd41; 
32'd550: dataIn2 = 32'd98; 
32'd551: dataIn2 = 32'd27; 
32'd552: dataIn2 = 32'd98; 
32'd553: dataIn2 = 32'd6; 
32'd554: dataIn2 = 32'd69; 
32'd555: dataIn2 = 32'd83; 
32'd556: dataIn2 = 32'd89; 
32'd557: dataIn2 = 32'd35; 
32'd558: dataIn2 = 32'd80; 
32'd559: dataIn2 = 32'd87; 
32'd560: dataIn2 = 32'd28; 
32'd561: dataIn2 = 32'd9; 
32'd562: dataIn2 = 32'd84; 
32'd563: dataIn2 = 32'd86; 
32'd564: dataIn2 = 32'd12; 
32'd565: dataIn2 = 32'd37; 
32'd566: dataIn2 = 32'd49; 
32'd567: dataIn2 = 32'd92; 
32'd568: dataIn2 = 32'd39; 
32'd569: dataIn2 = 32'd19; 
32'd570: dataIn2 = 32'd31; 
32'd571: dataIn2 = 32'd60; 
32'd572: dataIn2 = 32'd76; 
32'd573: dataIn2 = 32'd57; 
32'd574: dataIn2 = 32'd2; 
32'd575: dataIn2 = 32'd23; 
32'd576: dataIn2 = 32'd2; 
32'd577: dataIn2 = 32'd60; 
32'd578: dataIn2 = 32'd57; 
32'd579: dataIn2 = 32'd82; 
32'd580: dataIn2 = 32'd63; 
32'd581: dataIn2 = 32'd45; 
32'd582: dataIn2 = 32'd41; 
32'd583: dataIn2 = 32'd31; 
32'd584: dataIn2 = 32'd19; 
32'd585: dataIn2 = 32'd7; 
32'd586: dataIn2 = 32'd80; 
32'd587: dataIn2 = 32'd73; 
32'd588: dataIn2 = 32'd50; 
32'd589: dataIn2 = 32'd74; 
32'd590: dataIn2 = 32'd80; 
32'd591: dataIn2 = 32'd32; 
32'd592: dataIn2 = 32'd49; 
32'd593: dataIn2 = 32'd33; 
32'd594: dataIn2 = 32'd84; 
32'd595: dataIn2 = 32'd59; 
32'd596: dataIn2 = 32'd57; 
32'd597: dataIn2 = 32'd7; 
32'd598: dataIn2 = 32'd20; 
32'd599: dataIn2 = 32'd49; 
32'd600: dataIn2 = 32'd91; 
32'd601: dataIn2 = 32'd60; 
32'd602: dataIn2 = 32'd2; 
32'd603: dataIn2 = 32'd79; 
32'd604: dataIn2 = 32'd61; 
32'd605: dataIn2 = 32'd82; 
32'd606: dataIn2 = 32'd31; 
32'd607: dataIn2 = 32'd32; 
32'd608: dataIn2 = 32'd60; 
32'd609: dataIn2 = 32'd28; 
32'd610: dataIn2 = 32'd36; 
32'd611: dataIn2 = 32'd62; 
32'd612: dataIn2 = 32'd36; 
32'd613: dataIn2 = 32'd81; 
32'd614: dataIn2 = 32'd98; 
32'd615: dataIn2 = 32'd36; 
32'd616: dataIn2 = 32'd58; 
32'd617: dataIn2 = 32'd5; 
32'd618: dataIn2 = 32'd33; 
32'd619: dataIn2 = 32'd55; 
32'd620: dataIn2 = 32'd45; 
32'd621: dataIn2 = 32'd63; 
32'd622: dataIn2 = 32'd71; 
32'd623: dataIn2 = 32'd2; 
32'd624: dataIn2 = 32'd54; 
32'd625: dataIn2 = 32'd85; 
32'd626: dataIn2 = 32'd65; 
32'd627: dataIn2 = 32'd19; 
32'd628: dataIn2 = 32'd39; 
32'd629: dataIn2 = 32'd69; 
32'd630: dataIn2 = 32'd54; 
32'd631: dataIn2 = 32'd73; 
32'd632: dataIn2 = 32'd72; 
32'd633: dataIn2 = 32'd16; 
32'd634: dataIn2 = 32'd2; 
32'd635: dataIn2 = 32'd49; 
32'd636: dataIn2 = 32'd35; 
32'd637: dataIn2 = 32'd96; 
32'd638: dataIn2 = 32'd64; 
32'd639: dataIn2 = 32'd12; 
32'd640: dataIn2 = 32'd61; 
32'd641: dataIn2 = 32'd56; 
32'd642: dataIn2 = 32'd0; 
32'd643: dataIn2 = 32'd75; 
32'd644: dataIn2 = 32'd13; 
32'd645: dataIn2 = 32'd81; 
32'd646: dataIn2 = 32'd69; 
32'd647: dataIn2 = 32'd76; 
32'd648: dataIn2 = 32'd66; 
32'd649: dataIn2 = 32'd32; 
32'd650: dataIn2 = 32'd69; 
32'd651: dataIn2 = 32'd44; 
32'd652: dataIn2 = 32'd11; 
32'd653: dataIn2 = 32'd26; 
32'd654: dataIn2 = 32'd78; 
32'd655: dataIn2 = 32'd44; 
32'd656: dataIn2 = 32'd37; 
32'd657: dataIn2 = 32'd0; 
32'd658: dataIn2 = 32'd62; 
32'd659: dataIn2 = 32'd11; 
32'd660: dataIn2 = 32'd8; 
32'd661: dataIn2 = 32'd46; 
32'd662: dataIn2 = 32'd29; 
32'd663: dataIn2 = 32'd63; 
32'd664: dataIn2 = 32'd34; 
32'd665: dataIn2 = 32'd24; 
32'd666: dataIn2 = 32'd66; 
32'd667: dataIn2 = 32'd17; 
32'd668: dataIn2 = 32'd53; 
32'd669: dataIn2 = 32'd26; 
32'd670: dataIn2 = 32'd74; 
32'd671: dataIn2 = 32'd81; 
32'd672: dataIn2 = 32'd27; 
32'd673: dataIn2 = 32'd82; 
32'd674: dataIn2 = 32'd13; 
32'd675: dataIn2 = 32'd30; 
32'd676: dataIn2 = 32'd35; 
32'd677: dataIn2 = 32'd44; 
32'd678: dataIn2 = 32'd90; 
32'd679: dataIn2 = 32'd61; 
32'd680: dataIn2 = 32'd29; 
32'd681: dataIn2 = 32'd14; 
32'd682: dataIn2 = 32'd68; 
32'd683: dataIn2 = 32'd91; 
32'd684: dataIn2 = 32'd95; 
32'd685: dataIn2 = 32'd46; 
32'd686: dataIn2 = 32'd52; 
32'd687: dataIn2 = 32'd27; 
32'd688: dataIn2 = 32'd53; 
32'd689: dataIn2 = 32'd83; 
32'd690: dataIn2 = 32'd94; 
32'd691: dataIn2 = 32'd75; 
32'd692: dataIn2 = 32'd4; 
32'd693: dataIn2 = 32'd1; 
32'd694: dataIn2 = 32'd55; 
32'd695: dataIn2 = 32'd99; 
32'd696: dataIn2 = 32'd89; 
32'd697: dataIn2 = 32'd42; 
32'd698: dataIn2 = 32'd92; 
32'd699: dataIn2 = 32'd9; 
32'd700: dataIn2 = 32'd45; 
32'd701: dataIn2 = 32'd15; 
32'd702: dataIn2 = 32'd50; 
32'd703: dataIn2 = 32'd67; 
32'd704: dataIn2 = 32'd92; 
32'd705: dataIn2 = 32'd67; 
32'd706: dataIn2 = 32'd0; 
32'd707: dataIn2 = 32'd84; 
32'd708: dataIn2 = 32'd1; 
32'd709: dataIn2 = 32'd14; 
32'd710: dataIn2 = 32'd95; 
32'd711: dataIn2 = 32'd69; 
32'd712: dataIn2 = 32'd98; 
32'd713: dataIn2 = 32'd7; 
32'd714: dataIn2 = 32'd82; 
32'd715: dataIn2 = 32'd36; 
32'd716: dataIn2 = 32'd39; 
32'd717: dataIn2 = 32'd27; 
32'd718: dataIn2 = 32'd25; 
32'd719: dataIn2 = 32'd32; 
32'd720: dataIn2 = 32'd80; 
32'd721: dataIn2 = 32'd27; 
32'd722: dataIn2 = 32'd58; 
32'd723: dataIn2 = 32'd29; 
32'd724: dataIn2 = 32'd35; 
32'd725: dataIn2 = 32'd33; 
32'd726: dataIn2 = 32'd52; 
32'd727: dataIn2 = 32'd75; 
32'd728: dataIn2 = 32'd70; 
32'd729: dataIn2 = 32'd76; 
32'd730: dataIn2 = 32'd6; 
32'd731: dataIn2 = 32'd50; 
32'd732: dataIn2 = 32'd48; 
32'd733: dataIn2 = 32'd50; 
32'd734: dataIn2 = 32'd25; 
32'd735: dataIn2 = 32'd89; 
32'd736: dataIn2 = 32'd81; 
32'd737: dataIn2 = 32'd47; 
32'd738: dataIn2 = 32'd47; 
32'd739: dataIn2 = 32'd74; 
32'd740: dataIn2 = 32'd91; 
32'd741: dataIn2 = 32'd79; 
32'd742: dataIn2 = 32'd57; 
32'd743: dataIn2 = 32'd51; 
32'd744: dataIn2 = 32'd46; 
32'd745: dataIn2 = 32'd57; 
32'd746: dataIn2 = 32'd10; 
32'd747: dataIn2 = 32'd13; 
32'd748: dataIn2 = 32'd12; 
32'd749: dataIn2 = 32'd47; 
32'd750: dataIn2 = 32'd89; 
32'd751: dataIn2 = 32'd29; 
32'd752: dataIn2 = 32'd88; 
32'd753: dataIn2 = 32'd0; 
32'd754: dataIn2 = 32'd6; 
32'd755: dataIn2 = 32'd100; 
32'd756: dataIn2 = 32'd52; 
32'd757: dataIn2 = 32'd39; 
32'd758: dataIn2 = 32'd48; 
32'd759: dataIn2 = 32'd18; 
32'd760: dataIn2 = 32'd79; 
32'd761: dataIn2 = 32'd25; 
32'd762: dataIn2 = 32'd60; 
32'd763: dataIn2 = 32'd4; 
32'd764: dataIn2 = 32'd59; 
32'd765: dataIn2 = 32'd8; 
32'd766: dataIn2 = 32'd81; 
32'd767: dataIn2 = 32'd78; 
32'd768: dataIn2 = 32'd40; 
32'd769: dataIn2 = 32'd45; 
32'd770: dataIn2 = 32'd38; 
32'd771: dataIn2 = 32'd64; 
32'd772: dataIn2 = 32'd15; 
32'd773: dataIn2 = 32'd59; 
32'd774: dataIn2 = 32'd64; 
32'd775: dataIn2 = 32'd84; 
32'd776: dataIn2 = 32'd0; 
32'd777: dataIn2 = 32'd47; 
32'd778: dataIn2 = 32'd25; 
32'd779: dataIn2 = 32'd98; 
32'd780: dataIn2 = 32'd25; 
32'd781: dataIn2 = 32'd62; 
32'd782: dataIn2 = 32'd8; 
32'd783: dataIn2 = 32'd99; 
32'd784: dataIn2 = 32'd89; 
32'd785: dataIn2 = 32'd99; 
32'd786: dataIn2 = 32'd83; 
32'd787: dataIn2 = 32'd27; 
32'd788: dataIn2 = 32'd12; 
32'd789: dataIn2 = 32'd9; 
32'd790: dataIn2 = 32'd47; 
32'd791: dataIn2 = 32'd97; 
32'd792: dataIn2 = 32'd16; 
32'd793: dataIn2 = 32'd85; 
32'd794: dataIn2 = 32'd10; 
32'd795: dataIn2 = 32'd3; 
32'd796: dataIn2 = 32'd62; 
32'd797: dataIn2 = 32'd35; 
32'd798: dataIn2 = 32'd79; 
32'd799: dataIn2 = 32'd79; 
32'd800: dataIn2 = 32'd76; 
32'd801: dataIn2 = 32'd18; 
32'd802: dataIn2 = 32'd19; 
32'd803: dataIn2 = 32'd77; 
32'd804: dataIn2 = 32'd30; 
32'd805: dataIn2 = 32'd67; 
32'd806: dataIn2 = 32'd48; 
32'd807: dataIn2 = 32'd100; 
32'd808: dataIn2 = 32'd13; 
32'd809: dataIn2 = 32'd7; 
32'd810: dataIn2 = 32'd16; 
32'd811: dataIn2 = 32'd81; 
32'd812: dataIn2 = 32'd45; 
32'd813: dataIn2 = 32'd15; 
32'd814: dataIn2 = 32'd25; 
32'd815: dataIn2 = 32'd81; 
32'd816: dataIn2 = 32'd67; 
32'd817: dataIn2 = 32'd23; 
32'd818: dataIn2 = 32'd100; 
32'd819: dataIn2 = 32'd25; 
32'd820: dataIn2 = 32'd90; 
32'd821: dataIn2 = 32'd59; 
32'd822: dataIn2 = 32'd54; 
32'd823: dataIn2 = 32'd73; 
32'd824: dataIn2 = 32'd82; 
32'd825: dataIn2 = 32'd33; 
32'd826: dataIn2 = 32'd85; 
32'd827: dataIn2 = 32'd32; 
32'd828: dataIn2 = 32'd33; 
32'd829: dataIn2 = 32'd84; 
32'd830: dataIn2 = 32'd44; 
32'd831: dataIn2 = 32'd52; 
32'd832: dataIn2 = 32'd48; 
32'd833: dataIn2 = 32'd74; 
32'd834: dataIn2 = 32'd58; 
32'd835: dataIn2 = 32'd13; 
32'd836: dataIn2 = 32'd39; 
32'd837: dataIn2 = 32'd37; 
32'd838: dataIn2 = 32'd67; 
32'd839: dataIn2 = 32'd25; 
32'd840: dataIn2 = 32'd46; 
32'd841: dataIn2 = 32'd60; 
32'd842: dataIn2 = 32'd29; 
32'd843: dataIn2 = 32'd78; 
32'd844: dataIn2 = 32'd91; 
32'd845: dataIn2 = 32'd73; 
32'd846: dataIn2 = 32'd34; 
32'd847: dataIn2 = 32'd66; 
32'd848: dataIn2 = 32'd92; 
32'd849: dataIn2 = 32'd4; 
32'd850: dataIn2 = 32'd98; 
32'd851: dataIn2 = 32'd26; 
32'd852: dataIn2 = 32'd81; 
32'd853: dataIn2 = 32'd58; 
32'd854: dataIn2 = 32'd20; 
32'd855: dataIn2 = 32'd65; 
32'd856: dataIn2 = 32'd19; 
32'd857: dataIn2 = 32'd43; 
32'd858: dataIn2 = 32'd31; 
32'd859: dataIn2 = 32'd24; 
32'd860: dataIn2 = 32'd67; 
32'd861: dataIn2 = 32'd24; 
32'd862: dataIn2 = 32'd36; 
32'd863: dataIn2 = 32'd1; 
32'd864: dataIn2 = 32'd51; 
32'd865: dataIn2 = 32'd33; 
32'd866: dataIn2 = 32'd5; 
32'd867: dataIn2 = 32'd84; 
32'd868: dataIn2 = 32'd13; 
32'd869: dataIn2 = 32'd9; 
32'd870: dataIn2 = 32'd40; 
32'd871: dataIn2 = 32'd18; 
32'd872: dataIn2 = 32'd37; 
32'd873: dataIn2 = 32'd49; 
32'd874: dataIn2 = 32'd36; 
32'd875: dataIn2 = 32'd37; 
32'd876: dataIn2 = 32'd53; 
32'd877: dataIn2 = 32'd86; 
32'd878: dataIn2 = 32'd50; 
32'd879: dataIn2 = 32'd81; 
32'd880: dataIn2 = 32'd17; 
32'd881: dataIn2 = 32'd99; 
32'd882: dataIn2 = 32'd63; 
32'd883: dataIn2 = 32'd95; 
32'd884: dataIn2 = 32'd20; 
32'd885: dataIn2 = 32'd47; 
32'd886: dataIn2 = 32'd5; 
32'd887: dataIn2 = 32'd39; 
32'd888: dataIn2 = 32'd26; 
32'd889: dataIn2 = 32'd11; 
32'd890: dataIn2 = 32'd41; 
32'd891: dataIn2 = 32'd90; 
32'd892: dataIn2 = 32'd71; 
32'd893: dataIn2 = 32'd58; 
32'd894: dataIn2 = 32'd64; 
32'd895: dataIn2 = 32'd1; 
32'd896: dataIn2 = 32'd39; 
32'd897: dataIn2 = 32'd81; 
32'd898: dataIn2 = 32'd77; 
32'd899: dataIn2 = 32'd53; 
32'd900: dataIn2 = 32'd70; 
32'd901: dataIn2 = 32'd8; 
32'd902: dataIn2 = 32'd22; 
32'd903: dataIn2 = 32'd60; 
32'd904: dataIn2 = 32'd56; 
32'd905: dataIn2 = 32'd60; 
32'd906: dataIn2 = 32'd37; 
32'd907: dataIn2 = 32'd29; 
32'd908: dataIn2 = 32'd100; 
32'd909: dataIn2 = 32'd100; 
32'd910: dataIn2 = 32'd68; 
32'd911: dataIn2 = 32'd75; 
32'd912: dataIn2 = 32'd74; 
32'd913: dataIn2 = 32'd54; 
32'd914: dataIn2 = 32'd42; 
32'd915: dataIn2 = 32'd43; 
32'd916: dataIn2 = 32'd66; 
32'd917: dataIn2 = 32'd2; 
32'd918: dataIn2 = 32'd44; 
32'd919: dataIn2 = 32'd78; 
32'd920: dataIn2 = 32'd21; 
32'd921: dataIn2 = 32'd96; 
32'd922: dataIn2 = 32'd46; 
32'd923: dataIn2 = 32'd90; 
32'd924: dataIn2 = 32'd37; 
32'd925: dataIn2 = 32'd70; 
32'd926: dataIn2 = 32'd63; 
32'd927: dataIn2 = 32'd43; 
32'd928: dataIn2 = 32'd44; 
32'd929: dataIn2 = 32'd76; 
32'd930: dataIn2 = 32'd52; 
32'd931: dataIn2 = 32'd52; 
32'd932: dataIn2 = 32'd19; 
32'd933: dataIn2 = 32'd41; 
32'd934: dataIn2 = 32'd71; 
32'd935: dataIn2 = 32'd10; 
32'd936: dataIn2 = 32'd93; 
32'd937: dataIn2 = 32'd47; 
32'd938: dataIn2 = 32'd24; 
32'd939: dataIn2 = 32'd24; 
32'd940: dataIn2 = 32'd58; 
32'd941: dataIn2 = 32'd93; 
32'd942: dataIn2 = 32'd18; 
32'd943: dataIn2 = 32'd92; 
32'd944: dataIn2 = 32'd64; 
32'd945: dataIn2 = 32'd91; 
32'd946: dataIn2 = 32'd46; 
32'd947: dataIn2 = 32'd80; 
32'd948: dataIn2 = 32'd75; 
32'd949: dataIn2 = 32'd53; 
32'd950: dataIn2 = 32'd59; 
32'd951: dataIn2 = 32'd63; 
32'd952: dataIn2 = 32'd4; 
32'd953: dataIn2 = 32'd19; 
32'd954: dataIn2 = 32'd48; 
32'd955: dataIn2 = 32'd36; 
32'd956: dataIn2 = 32'd71; 
32'd957: dataIn2 = 32'd43; 
32'd958: dataIn2 = 32'd22; 
32'd959: dataIn2 = 32'd48; 
32'd960: dataIn2 = 32'd76; 
32'd961: dataIn2 = 32'd85; 
32'd962: dataIn2 = 32'd24; 
32'd963: dataIn2 = 32'd37; 
32'd964: dataIn2 = 32'd53; 
32'd965: dataIn2 = 32'd43; 
32'd966: dataIn2 = 32'd95; 
32'd967: dataIn2 = 32'd16; 
32'd968: dataIn2 = 32'd2; 
32'd969: dataIn2 = 32'd29; 
32'd970: dataIn2 = 32'd38; 
32'd971: dataIn2 = 32'd69; 
32'd972: dataIn2 = 32'd54; 
32'd973: dataIn2 = 32'd12; 
32'd974: dataIn2 = 32'd49; 
32'd975: dataIn2 = 32'd40; 
32'd976: dataIn2 = 32'd75; 
32'd977: dataIn2 = 32'd96; 
32'd978: dataIn2 = 32'd48; 
32'd979: dataIn2 = 32'd65; 
32'd980: dataIn2 = 32'd82; 
32'd981: dataIn2 = 32'd56; 
32'd982: dataIn2 = 32'd55; 
32'd983: dataIn2 = 32'd69; 
32'd984: dataIn2 = 32'd12; 
32'd985: dataIn2 = 32'd75; 
32'd986: dataIn2 = 32'd24; 
32'd987: dataIn2 = 32'd11; 
32'd988: dataIn2 = 32'd50; 
32'd989: dataIn2 = 32'd44; 
32'd990: dataIn2 = 32'd88; 
32'd991: dataIn2 = 32'd56; 
32'd992: dataIn2 = 32'd90; 
32'd993: dataIn2 = 32'd72; 
32'd994: dataIn2 = 32'd6; 
32'd995: dataIn2 = 32'd76; 
32'd996: dataIn2 = 32'd7; 
32'd997: dataIn2 = 32'd80; 
32'd998: dataIn2 = 32'd93; 
32'd999: dataIn2 = 32'd18; 
32'd1000: dataIn2 = 32'd30; 
32'd1001: dataIn2 = 32'd89; 
32'd1002: dataIn2 = 32'd52; 
32'd1003: dataIn2 = 32'd31; 
32'd1004: dataIn2 = 32'd12; 
32'd1005: dataIn2 = 32'd60; 
32'd1006: dataIn2 = 32'd22; 
32'd1007: dataIn2 = 32'd13; 
32'd1008: dataIn2 = 32'd75; 
32'd1009: dataIn2 = 32'd5; 
32'd1010: dataIn2 = 32'd11; 
32'd1011: dataIn2 = 32'd78; 
32'd1012: dataIn2 = 32'd6; 
32'd1013: dataIn2 = 32'd69; 
32'd1014: dataIn2 = 32'd50; 
32'd1015: dataIn2 = 32'd21; 
32'd1016: dataIn2 = 32'd77; 
32'd1017: dataIn2 = 32'd67; 
32'd1018: dataIn2 = 32'd98; 
32'd1019: dataIn2 = 32'd88; 
32'd1020: dataIn2 = 32'd24; 
32'd1021: dataIn2 = 32'd79; 
32'd1022: dataIn2 = 32'd0; 
32'd1023: dataIn2 = 32'd30; 
32'd1024: dataIn2 = 32'd47; 
32'd1025: dataIn2 = 32'd71; 
32'd1026: dataIn2 = 32'd65; 
32'd1027: dataIn2 = 32'd52; 
32'd1028: dataIn2 = 32'd13; 
32'd1029: dataIn2 = 32'd57; 
32'd1030: dataIn2 = 32'd76; 
32'd1031: dataIn2 = 32'd54; 
32'd1032: dataIn2 = 32'd37; 
32'd1033: dataIn2 = 32'd21; 
32'd1034: dataIn2 = 32'd77; 
32'd1035: dataIn2 = 32'd79; 
32'd1036: dataIn2 = 32'd25; 
32'd1037: dataIn2 = 32'd51; 
32'd1038: dataIn2 = 32'd17; 
32'd1039: dataIn2 = 32'd71; 
32'd1040: dataIn2 = 32'd23; 
32'd1041: dataIn2 = 32'd17; 
32'd1042: dataIn2 = 32'd91; 
32'd1043: dataIn2 = 32'd67; 
32'd1044: dataIn2 = 32'd7; 
32'd1045: dataIn2 = 32'd31; 
32'd1046: dataIn2 = 32'd69; 
32'd1047: dataIn2 = 32'd96; 
32'd1048: dataIn2 = 32'd40; 
32'd1049: dataIn2 = 32'd81; 
32'd1050: dataIn2 = 32'd84; 
32'd1051: dataIn2 = 32'd26; 
32'd1052: dataIn2 = 32'd18; 
32'd1053: dataIn2 = 32'd37; 
32'd1054: dataIn2 = 32'd43; 
32'd1055: dataIn2 = 32'd64; 
32'd1056: dataIn2 = 32'd17; 
32'd1057: dataIn2 = 32'd80; 
32'd1058: dataIn2 = 32'd46; 
32'd1059: dataIn2 = 32'd49; 
32'd1060: dataIn2 = 32'd8; 
32'd1061: dataIn2 = 32'd47; 
32'd1062: dataIn2 = 32'd87; 
32'd1063: dataIn2 = 32'd1; 
32'd1064: dataIn2 = 32'd96; 
32'd1065: dataIn2 = 32'd47; 
32'd1066: dataIn2 = 32'd11; 
32'd1067: dataIn2 = 32'd14; 
32'd1068: dataIn2 = 32'd3; 
32'd1069: dataIn2 = 32'd10; 
32'd1070: dataIn2 = 32'd80; 
32'd1071: dataIn2 = 32'd52; 
32'd1072: dataIn2 = 32'd99; 
32'd1073: dataIn2 = 32'd92; 
32'd1074: dataIn2 = 32'd64; 
32'd1075: dataIn2 = 32'd42; 
32'd1076: dataIn2 = 32'd6; 
32'd1077: dataIn2 = 32'd98; 
32'd1078: dataIn2 = 32'd63; 
32'd1079: dataIn2 = 32'd82; 
32'd1080: dataIn2 = 32'd14; 
32'd1081: dataIn2 = 32'd9; 
32'd1082: dataIn2 = 32'd91; 
32'd1083: dataIn2 = 32'd35; 
32'd1084: dataIn2 = 32'd50; 
32'd1085: dataIn2 = 32'd76; 
32'd1086: dataIn2 = 32'd11; 
32'd1087: dataIn2 = 32'd65; 
32'd1088: dataIn2 = 32'd3; 
32'd1089: dataIn2 = 32'd83; 
32'd1090: dataIn2 = 32'd79; 
32'd1091: dataIn2 = 32'd31; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_new_32_10.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
