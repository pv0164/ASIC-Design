//64x64 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 2048 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,addr1,addr2,dataIn1,dataIn2,Rst,csize,RD);  
//frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  wdata_col_base = 32'd660 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #41140; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd660: dataIn1 = 32'd37; 
32'd661: dataIn1 = 32'd5; 
32'd662: dataIn1 = 32'd41; 
32'd663: dataIn1 = 32'd62; 
32'd664: dataIn1 = 32'd52; 
32'd665: dataIn1 = 32'd13; 
32'd666: dataIn1 = 32'd32; 
32'd667: dataIn1 = 32'd40; 
32'd668: dataIn1 = 32'd5; 
32'd669: dataIn1 = 32'd15; 
32'd670: dataIn1 = 32'd11; 
32'd671: dataIn1 = 32'd10; 
32'd672: dataIn1 = 32'd19; 
32'd673: dataIn1 = 32'd45; 
32'd674: dataIn1 = 32'd54; 
32'd675: dataIn1 = 32'd63; 
32'd676: dataIn1 = 32'd49; 
32'd677: dataIn1 = 32'd57; 
32'd678: dataIn1 = 32'd52; 
32'd679: dataIn1 = 32'd57; 
32'd680: dataIn1 = 32'd16; 
32'd681: dataIn1 = 32'd0; 
32'd682: dataIn1 = 32'd13; 
32'd683: dataIn1 = 32'd43; 
32'd684: dataIn1 = 32'd36; 
32'd685: dataIn1 = 32'd48; 
32'd686: dataIn1 = 32'd10; 
32'd687: dataIn1 = 32'd36; 
32'd688: dataIn1 = 32'd44; 
32'd689: dataIn1 = 32'd9; 
32'd690: dataIn1 = 32'd39; 
32'd691: dataIn1 = 32'd41; 
32'd692: dataIn1 = 32'd26; 
32'd693: dataIn1 = 32'd19; 
32'd694: dataIn1 = 32'd52; 
32'd695: dataIn1 = 32'd62; 
32'd696: dataIn1 = 32'd24; 
32'd697: dataIn1 = 32'd53; 
32'd698: dataIn1 = 32'd62; 
32'd699: dataIn1 = 32'd13; 
32'd700: dataIn1 = 32'd55; 
32'd701: dataIn1 = 32'd17; 
32'd702: dataIn1 = 32'd17; 
32'd703: dataIn1 = 32'd27; 
32'd704: dataIn1 = 32'd55; 
32'd705: dataIn1 = 32'd32; 
32'd706: dataIn1 = 32'd49; 
32'd707: dataIn1 = 32'd58; 
32'd708: dataIn1 = 32'd57; 
32'd709: dataIn1 = 32'd12; 
32'd710: dataIn1 = 32'd48; 
32'd711: dataIn1 = 32'd30; 
32'd712: dataIn1 = 32'd20; 
32'd713: dataIn1 = 32'd36; 
32'd714: dataIn1 = 32'd30; 
32'd715: dataIn1 = 32'd14; 
32'd716: dataIn1 = 32'd5; 
32'd717: dataIn1 = 32'd29; 
32'd718: dataIn1 = 32'd62; 
32'd719: dataIn1 = 32'd22; 
32'd720: dataIn1 = 32'd6; 
32'd721: dataIn1 = 32'd14; 
32'd722: dataIn1 = 32'd7; 
32'd723: dataIn1 = 32'd37; 
32'd724: dataIn1 = 32'd17; 
32'd725: dataIn1 = 32'd51; 
32'd726: dataIn1 = 32'd50; 
32'd727: dataIn1 = 32'd9; 
32'd728: dataIn1 = 32'd12; 
32'd729: dataIn1 = 32'd23; 
32'd730: dataIn1 = 32'd2; 
32'd731: dataIn1 = 32'd1; 
32'd732: dataIn1 = 32'd54; 
32'd733: dataIn1 = 32'd43; 
32'd734: dataIn1 = 32'd3; 
32'd735: dataIn1 = 32'd55; 
32'd736: dataIn1 = 32'd0; 
32'd737: dataIn1 = 32'd16; 
32'd738: dataIn1 = 32'd22; 
32'd739: dataIn1 = 32'd42; 
32'd740: dataIn1 = 32'd27; 
32'd741: dataIn1 = 32'd57; 
32'd742: dataIn1 = 32'd55; 
32'd743: dataIn1 = 32'd6; 
32'd744: dataIn1 = 32'd42; 
32'd745: dataIn1 = 32'd1; 
32'd746: dataIn1 = 32'd35; 
32'd747: dataIn1 = 32'd46; 
32'd748: dataIn1 = 32'd28; 
32'd749: dataIn1 = 32'd7; 
32'd750: dataIn1 = 32'd26; 
32'd751: dataIn1 = 32'd62; 
32'd752: dataIn1 = 32'd19; 
32'd753: dataIn1 = 32'd48; 
32'd754: dataIn1 = 32'd26; 
32'd755: dataIn1 = 32'd8; 
32'd756: dataIn1 = 32'd30; 
32'd757: dataIn1 = 32'd8; 
32'd758: dataIn1 = 32'd43; 
32'd759: dataIn1 = 32'd48; 
32'd760: dataIn1 = 32'd51; 
32'd761: dataIn1 = 32'd6; 
32'd762: dataIn1 = 32'd44; 
32'd763: dataIn1 = 32'd21; 
32'd764: dataIn1 = 32'd24; 
32'd765: dataIn1 = 32'd8; 
32'd766: dataIn1 = 32'd52; 
32'd767: dataIn1 = 32'd46; 
32'd768: dataIn1 = 32'd26; 
32'd769: dataIn1 = 32'd63; 
32'd770: dataIn1 = 32'd32; 
32'd771: dataIn1 = 32'd1; 
32'd772: dataIn1 = 32'd57; 
32'd773: dataIn1 = 32'd42; 
32'd774: dataIn1 = 32'd14; 
32'd775: dataIn1 = 32'd38; 
32'd776: dataIn1 = 32'd34; 
32'd777: dataIn1 = 32'd37; 
32'd778: dataIn1 = 32'd2; 
32'd779: dataIn1 = 32'd31; 
32'd780: dataIn1 = 32'd36; 
32'd781: dataIn1 = 32'd33; 
32'd782: dataIn1 = 32'd17; 
32'd783: dataIn1 = 32'd47; 
32'd784: dataIn1 = 32'd0; 
32'd785: dataIn1 = 32'd27; 
32'd786: dataIn1 = 32'd34; 
32'd787: dataIn1 = 32'd35; 
32'd788: dataIn1 = 32'd19; 
32'd789: dataIn1 = 32'd50; 
32'd790: dataIn1 = 32'd43; 
32'd791: dataIn1 = 32'd42; 
32'd792: dataIn1 = 32'd62; 
32'd793: dataIn1 = 32'd24; 
32'd794: dataIn1 = 32'd41; 
32'd795: dataIn1 = 32'd59; 
32'd796: dataIn1 = 32'd32; 
32'd797: dataIn1 = 32'd11; 
32'd798: dataIn1 = 32'd29; 
32'd799: dataIn1 = 32'd55; 
32'd800: dataIn1 = 32'd37; 
32'd801: dataIn1 = 32'd38; 
32'd802: dataIn1 = 32'd50; 
32'd803: dataIn1 = 32'd33; 
32'd804: dataIn1 = 32'd49; 
32'd805: dataIn1 = 32'd26; 
32'd806: dataIn1 = 32'd40; 
32'd807: dataIn1 = 32'd44; 
32'd808: dataIn1 = 32'd23; 
32'd809: dataIn1 = 32'd59; 
32'd810: dataIn1 = 32'd47; 
32'd811: dataIn1 = 32'd17; 
32'd812: dataIn1 = 32'd51; 
32'd813: dataIn1 = 32'd61; 
32'd814: dataIn1 = 32'd29; 
32'd815: dataIn1 = 32'd59; 
32'd816: dataIn1 = 32'd4; 
32'd817: dataIn1 = 32'd12; 
32'd818: dataIn1 = 32'd7; 
32'd819: dataIn1 = 32'd55; 
32'd820: dataIn1 = 32'd56; 
32'd821: dataIn1 = 32'd15; 
32'd822: dataIn1 = 32'd17; 
32'd823: dataIn1 = 32'd23; 
32'd824: dataIn1 = 32'd7; 
32'd825: dataIn1 = 32'd57; 
32'd826: dataIn1 = 32'd57; 
32'd827: dataIn1 = 32'd56; 
32'd828: dataIn1 = 32'd62; 
32'd829: dataIn1 = 32'd38; 
32'd830: dataIn1 = 32'd44; 
32'd831: dataIn1 = 32'd24; 
32'd832: dataIn1 = 32'd14; 
32'd833: dataIn1 = 32'd10; 
32'd834: dataIn1 = 32'd61; 
32'd835: dataIn1 = 32'd30; 
32'd836: dataIn1 = 32'd40; 
32'd837: dataIn1 = 32'd59; 
32'd838: dataIn1 = 32'd37; 
32'd839: dataIn1 = 32'd30; 
32'd840: dataIn1 = 32'd26; 
32'd841: dataIn1 = 32'd43; 
32'd842: dataIn1 = 32'd0; 
32'd843: dataIn1 = 32'd39; 
32'd844: dataIn1 = 32'd59; 
32'd845: dataIn1 = 32'd44; 
32'd846: dataIn1 = 32'd42; 
32'd847: dataIn1 = 32'd21; 
32'd848: dataIn1 = 32'd4; 
32'd849: dataIn1 = 32'd27; 
32'd850: dataIn1 = 32'd19; 
32'd851: dataIn1 = 32'd59; 
32'd852: dataIn1 = 32'd8; 
32'd853: dataIn1 = 32'd63; 
32'd854: dataIn1 = 32'd22; 
32'd855: dataIn1 = 32'd33; 
32'd856: dataIn1 = 32'd63; 
32'd857: dataIn1 = 32'd47; 
32'd858: dataIn1 = 32'd44; 
32'd859: dataIn1 = 32'd17; 
32'd860: dataIn1 = 32'd55; 
32'd861: dataIn1 = 32'd41; 
32'd862: dataIn1 = 32'd58; 
32'd863: dataIn1 = 32'd23; 
32'd864: dataIn1 = 32'd6; 
32'd865: dataIn1 = 32'd59; 
32'd866: dataIn1 = 32'd8; 
32'd867: dataIn1 = 32'd23; 
32'd868: dataIn1 = 32'd25; 
32'd869: dataIn1 = 32'd15; 
32'd870: dataIn1 = 32'd21; 
32'd871: dataIn1 = 32'd56; 
32'd872: dataIn1 = 32'd15; 
32'd873: dataIn1 = 32'd52; 
32'd874: dataIn1 = 32'd60; 
32'd875: dataIn1 = 32'd14; 
32'd876: dataIn1 = 32'd53; 
32'd877: dataIn1 = 32'd22; 
32'd878: dataIn1 = 32'd15; 
32'd879: dataIn1 = 32'd36; 
32'd880: dataIn1 = 32'd4; 
32'd881: dataIn1 = 32'd20; 
32'd882: dataIn1 = 32'd38; 
32'd883: dataIn1 = 32'd24; 
32'd884: dataIn1 = 32'd62; 
32'd885: dataIn1 = 32'd34; 
32'd886: dataIn1 = 32'd57; 
32'd887: dataIn1 = 32'd49; 
32'd888: dataIn1 = 32'd48; 
32'd889: dataIn1 = 32'd31; 
32'd890: dataIn1 = 32'd6; 
32'd891: dataIn1 = 32'd51; 
32'd892: dataIn1 = 32'd17; 
32'd893: dataIn1 = 32'd17; 
32'd894: dataIn1 = 32'd46; 
32'd895: dataIn1 = 32'd61; 
32'd896: dataIn1 = 32'd59; 
32'd897: dataIn1 = 32'd36; 
32'd898: dataIn1 = 32'd31; 
32'd899: dataIn1 = 32'd26; 
32'd900: dataIn1 = 32'd42; 
32'd901: dataIn1 = 32'd59; 
32'd902: dataIn1 = 32'd51; 
32'd903: dataIn1 = 32'd61; 
32'd904: dataIn1 = 32'd28; 
32'd905: dataIn1 = 32'd61; 
32'd906: dataIn1 = 32'd32; 
32'd907: dataIn1 = 32'd25; 
32'd908: dataIn1 = 32'd1; 
32'd909: dataIn1 = 32'd63; 
32'd910: dataIn1 = 32'd0; 
32'd911: dataIn1 = 32'd41; 
32'd912: dataIn1 = 32'd38; 
32'd913: dataIn1 = 32'd14; 
32'd914: dataIn1 = 32'd21; 
32'd915: dataIn1 = 32'd26; 
32'd916: dataIn1 = 32'd24; 
32'd917: dataIn1 = 32'd36; 
32'd918: dataIn1 = 32'd22; 
32'd919: dataIn1 = 32'd43; 
32'd920: dataIn1 = 32'd61; 
32'd921: dataIn1 = 32'd54; 
32'd922: dataIn1 = 32'd23; 
32'd923: dataIn1 = 32'd13; 
32'd924: dataIn1 = 32'd57; 
32'd925: dataIn1 = 32'd37; 
32'd926: dataIn1 = 32'd48; 
32'd927: dataIn1 = 32'd42; 
32'd928: dataIn1 = 32'd54; 
32'd929: dataIn1 = 32'd30; 
32'd930: dataIn1 = 32'd39; 
32'd931: dataIn1 = 32'd19; 
32'd932: dataIn1 = 32'd53; 
32'd933: dataIn1 = 32'd53; 
32'd934: dataIn1 = 32'd50; 
32'd935: dataIn1 = 32'd46; 
32'd936: dataIn1 = 32'd32; 
32'd937: dataIn1 = 32'd61; 
32'd938: dataIn1 = 32'd37; 
32'd939: dataIn1 = 32'd39; 
32'd940: dataIn1 = 32'd43; 
32'd941: dataIn1 = 32'd38; 
32'd942: dataIn1 = 32'd8; 
32'd943: dataIn1 = 32'd10; 
32'd944: dataIn1 = 32'd36; 
32'd945: dataIn1 = 32'd54; 
32'd946: dataIn1 = 32'd59; 
32'd947: dataIn1 = 32'd29; 
32'd948: dataIn1 = 32'd18; 
32'd949: dataIn1 = 32'd50; 
32'd950: dataIn1 = 32'd52; 
32'd951: dataIn1 = 32'd8; 
32'd952: dataIn1 = 32'd6; 
32'd953: dataIn1 = 32'd54; 
32'd954: dataIn1 = 32'd62; 
32'd955: dataIn1 = 32'd21; 
32'd956: dataIn1 = 32'd3; 
32'd957: dataIn1 = 32'd11; 
32'd958: dataIn1 = 32'd39; 
32'd959: dataIn1 = 32'd52; 
32'd960: dataIn1 = 32'd3; 
32'd961: dataIn1 = 32'd53; 
32'd962: dataIn1 = 32'd13; 
32'd963: dataIn1 = 32'd44; 
32'd964: dataIn1 = 32'd2; 
32'd965: dataIn1 = 32'd59; 
32'd966: dataIn1 = 32'd18; 
32'd967: dataIn1 = 32'd12; 
32'd968: dataIn1 = 32'd0; 
32'd969: dataIn1 = 32'd27; 
32'd970: dataIn1 = 32'd60; 
32'd971: dataIn1 = 32'd19; 
32'd972: dataIn1 = 32'd22; 
32'd973: dataIn1 = 32'd44; 
32'd974: dataIn1 = 32'd27; 
32'd975: dataIn1 = 32'd44; 
32'd976: dataIn1 = 32'd55; 
32'd977: dataIn1 = 32'd49; 
32'd978: dataIn1 = 32'd41; 
32'd979: dataIn1 = 32'd47; 
32'd980: dataIn1 = 32'd42; 
32'd981: dataIn1 = 32'd59; 
32'd982: dataIn1 = 32'd42; 
32'd983: dataIn1 = 32'd0; 
32'd984: dataIn1 = 32'd55; 
32'd985: dataIn1 = 32'd6; 
32'd986: dataIn1 = 32'd38; 
32'd987: dataIn1 = 32'd27; 
32'd988: dataIn1 = 32'd46; 
32'd989: dataIn1 = 32'd44; 
32'd990: dataIn1 = 32'd56; 
32'd991: dataIn1 = 32'd63; 
32'd992: dataIn1 = 32'd56; 
32'd993: dataIn1 = 32'd40; 
32'd994: dataIn1 = 32'd49; 
32'd995: dataIn1 = 32'd12; 
32'd996: dataIn1 = 32'd45; 
32'd997: dataIn1 = 32'd38; 
32'd998: dataIn1 = 32'd49; 
32'd999: dataIn1 = 32'd17; 
32'd1000: dataIn1 = 32'd59; 
32'd1001: dataIn1 = 32'd54; 
32'd1002: dataIn1 = 32'd57; 
32'd1003: dataIn1 = 32'd34; 
32'd1004: dataIn1 = 32'd39; 
32'd1005: dataIn1 = 32'd52; 
32'd1006: dataIn1 = 32'd4; 
32'd1007: dataIn1 = 32'd18; 
32'd1008: dataIn1 = 32'd17; 
32'd1009: dataIn1 = 32'd57; 
32'd1010: dataIn1 = 32'd59; 
32'd1011: dataIn1 = 32'd62; 
32'd1012: dataIn1 = 32'd12; 
32'd1013: dataIn1 = 32'd12; 
32'd1014: dataIn1 = 32'd20; 
32'd1015: dataIn1 = 32'd12; 
32'd1016: dataIn1 = 32'd8; 
32'd1017: dataIn1 = 32'd31; 
32'd1018: dataIn1 = 32'd27; 
32'd1019: dataIn1 = 32'd52; 
32'd1020: dataIn1 = 32'd28; 
32'd1021: dataIn1 = 32'd6; 
32'd1022: dataIn1 = 32'd39; 
32'd1023: dataIn1 = 32'd23; 
32'd1024: dataIn1 = 32'd18; 
32'd1025: dataIn1 = 32'd53; 
32'd1026: dataIn1 = 32'd61; 
32'd1027: dataIn1 = 32'd12; 
32'd1028: dataIn1 = 32'd56; 
32'd1029: dataIn1 = 32'd18; 
32'd1030: dataIn1 = 32'd25; 
32'd1031: dataIn1 = 32'd58; 
32'd1032: dataIn1 = 32'd35; 
32'd1033: dataIn1 = 32'd32; 
32'd1034: dataIn1 = 32'd21; 
32'd1035: dataIn1 = 32'd14; 
32'd1036: dataIn1 = 32'd23; 
32'd1037: dataIn1 = 32'd63; 
32'd1038: dataIn1 = 32'd1; 
32'd1039: dataIn1 = 32'd38; 
32'd1040: dataIn1 = 32'd43; 
32'd1041: dataIn1 = 32'd10; 
32'd1042: dataIn1 = 32'd45; 
32'd1043: dataIn1 = 32'd15; 
32'd1044: dataIn1 = 32'd38; 
32'd1045: dataIn1 = 32'd45; 
32'd1046: dataIn1 = 32'd10; 
32'd1047: dataIn1 = 32'd58; 
32'd1048: dataIn1 = 32'd28; 
32'd1049: dataIn1 = 32'd46; 
32'd1050: dataIn1 = 32'd39; 
32'd1051: dataIn1 = 32'd17; 
32'd1052: dataIn1 = 32'd23; 
32'd1053: dataIn1 = 32'd24; 
32'd1054: dataIn1 = 32'd25; 
32'd1055: dataIn1 = 32'd49; 
32'd1056: dataIn1 = 32'd29; 
32'd1057: dataIn1 = 32'd45; 
32'd1058: dataIn1 = 32'd10; 
32'd1059: dataIn1 = 32'd51; 
32'd1060: dataIn1 = 32'd8; 
32'd1061: dataIn1 = 32'd48; 
32'd1062: dataIn1 = 32'd52; 
32'd1063: dataIn1 = 32'd34; 
32'd1064: dataIn1 = 32'd33; 
32'd1065: dataIn1 = 32'd9; 
32'd1066: dataIn1 = 32'd19; 
32'd1067: dataIn1 = 32'd14; 
32'd1068: dataIn1 = 32'd10; 
32'd1069: dataIn1 = 32'd11; 
32'd1070: dataIn1 = 32'd42; 
32'd1071: dataIn1 = 32'd16; 
32'd1072: dataIn1 = 32'd43; 
32'd1073: dataIn1 = 32'd2; 
32'd1074: dataIn1 = 32'd38; 
32'd1075: dataIn1 = 32'd28; 
32'd1076: dataIn1 = 32'd4; 
32'd1077: dataIn1 = 32'd43; 
32'd1078: dataIn1 = 32'd40; 
32'd1079: dataIn1 = 32'd33; 
32'd1080: dataIn1 = 32'd48; 
32'd1081: dataIn1 = 32'd44; 
32'd1082: dataIn1 = 32'd23; 
32'd1083: dataIn1 = 32'd34; 
32'd1084: dataIn1 = 32'd2; 
32'd1085: dataIn1 = 32'd1; 
32'd1086: dataIn1 = 32'd1; 
32'd1087: dataIn1 = 32'd27; 
32'd1088: dataIn1 = 32'd24; 
32'd1089: dataIn1 = 32'd53; 
32'd1090: dataIn1 = 32'd20; 
32'd1091: dataIn1 = 32'd1; 
32'd1092: dataIn1 = 32'd7; 
32'd1093: dataIn1 = 32'd11; 
32'd1094: dataIn1 = 32'd15; 
32'd1095: dataIn1 = 32'd54; 
32'd1096: dataIn1 = 32'd35; 
32'd1097: dataIn1 = 32'd25; 
32'd1098: dataIn1 = 32'd45; 
32'd1099: dataIn1 = 32'd53; 
32'd1100: dataIn1 = 32'd12; 
32'd1101: dataIn1 = 32'd48; 
32'd1102: dataIn1 = 32'd56; 
32'd1103: dataIn1 = 32'd63; 
32'd1104: dataIn1 = 32'd54; 
32'd1105: dataIn1 = 32'd30; 
32'd1106: dataIn1 = 32'd26; 
32'd1107: dataIn1 = 32'd35; 
32'd1108: dataIn1 = 32'd45; 
32'd1109: dataIn1 = 32'd41; 
32'd1110: dataIn1 = 32'd55; 
32'd1111: dataIn1 = 32'd59; 
32'd1112: dataIn1 = 32'd4; 
32'd1113: dataIn1 = 32'd13; 
32'd1114: dataIn1 = 32'd18; 
32'd1115: dataIn1 = 32'd48; 
32'd1116: dataIn1 = 32'd45; 
32'd1117: dataIn1 = 32'd25; 
32'd1118: dataIn1 = 32'd13; 
32'd1119: dataIn1 = 32'd41; 
32'd1120: dataIn1 = 32'd20; 
32'd1121: dataIn1 = 32'd56; 
32'd1122: dataIn1 = 32'd41; 
32'd1123: dataIn1 = 32'd35; 
32'd1124: dataIn1 = 32'd39; 
32'd1125: dataIn1 = 32'd1; 
32'd1126: dataIn1 = 32'd8; 
32'd1127: dataIn1 = 32'd8; 
32'd1128: dataIn1 = 32'd12; 
32'd1129: dataIn1 = 32'd11; 
32'd1130: dataIn1 = 32'd57; 
32'd1131: dataIn1 = 32'd9; 
32'd1132: dataIn1 = 32'd21; 
32'd1133: dataIn1 = 32'd5; 
32'd1134: dataIn1 = 32'd45; 
32'd1135: dataIn1 = 32'd48; 
32'd1136: dataIn1 = 32'd44; 
32'd1137: dataIn1 = 32'd61; 
32'd1138: dataIn1 = 32'd57; 
32'd1139: dataIn1 = 32'd47; 
32'd1140: dataIn1 = 32'd43; 
32'd1141: dataIn1 = 32'd14; 
32'd1142: dataIn1 = 32'd45; 
32'd1143: dataIn1 = 32'd4; 
32'd1144: dataIn1 = 32'd41; 
32'd1145: dataIn1 = 32'd62; 
32'd1146: dataIn1 = 32'd26; 
32'd1147: dataIn1 = 32'd35; 
32'd1148: dataIn1 = 32'd25; 
32'd1149: dataIn1 = 32'd26; 
32'd1150: dataIn1 = 32'd45; 
32'd1151: dataIn1 = 32'd1; 
32'd1152: dataIn1 = 32'd38; 
32'd1153: dataIn1 = 32'd39; 
32'd1154: dataIn1 = 32'd8; 
32'd1155: dataIn1 = 32'd53; 
32'd1156: dataIn1 = 32'd52; 
32'd1157: dataIn1 = 32'd63; 
32'd1158: dataIn1 = 32'd59; 
32'd1159: dataIn1 = 32'd48; 
32'd1160: dataIn1 = 32'd55; 
32'd1161: dataIn1 = 32'd5; 
32'd1162: dataIn1 = 32'd12; 
32'd1163: dataIn1 = 32'd38; 
32'd1164: dataIn1 = 32'd20; 
32'd1165: dataIn1 = 32'd19; 
32'd1166: dataIn1 = 32'd58; 
32'd1167: dataIn1 = 32'd37; 
32'd1168: dataIn1 = 32'd34; 
32'd1169: dataIn1 = 32'd55; 
32'd1170: dataIn1 = 32'd36; 
32'd1171: dataIn1 = 32'd17; 
32'd1172: dataIn1 = 32'd45; 
32'd1173: dataIn1 = 32'd18; 
32'd1174: dataIn1 = 32'd35; 
32'd1175: dataIn1 = 32'd25; 
32'd1176: dataIn1 = 32'd47; 
32'd1177: dataIn1 = 32'd57; 
32'd1178: dataIn1 = 32'd44; 
32'd1179: dataIn1 = 32'd2; 
32'd1180: dataIn1 = 32'd20; 
32'd1181: dataIn1 = 32'd16; 
32'd1182: dataIn1 = 32'd2; 
32'd1183: dataIn1 = 32'd28; 
32'd1184: dataIn1 = 32'd6; 
32'd1185: dataIn1 = 32'd46; 
32'd1186: dataIn1 = 32'd14; 
32'd1187: dataIn1 = 32'd29; 
32'd1188: dataIn1 = 32'd63; 
32'd1189: dataIn1 = 32'd59; 
32'd1190: dataIn1 = 32'd59; 
32'd1191: dataIn1 = 32'd55; 
32'd1192: dataIn1 = 32'd36; 
32'd1193: dataIn1 = 32'd7; 
32'd1194: dataIn1 = 32'd62; 
32'd1195: dataIn1 = 32'd21; 
32'd1196: dataIn1 = 32'd50; 
32'd1197: dataIn1 = 32'd54; 
32'd1198: dataIn1 = 32'd5; 
32'd1199: dataIn1 = 32'd6; 
32'd1200: dataIn1 = 32'd2; 
32'd1201: dataIn1 = 32'd25; 
32'd1202: dataIn1 = 32'd24; 
32'd1203: dataIn1 = 32'd42; 
32'd1204: dataIn1 = 32'd52; 
32'd1205: dataIn1 = 32'd56; 
32'd1206: dataIn1 = 32'd38; 
32'd1207: dataIn1 = 32'd51; 
32'd1208: dataIn1 = 32'd61; 
32'd1209: dataIn1 = 32'd34; 
32'd1210: dataIn1 = 32'd59; 
32'd1211: dataIn1 = 32'd54; 
32'd1212: dataIn1 = 32'd10; 
32'd1213: dataIn1 = 32'd33; 
32'd1214: dataIn1 = 32'd27; 
32'd1215: dataIn1 = 32'd37; 
32'd1216: dataIn1 = 32'd26; 
32'd1217: dataIn1 = 32'd39; 
32'd1218: dataIn1 = 32'd59; 
32'd1219: dataIn1 = 32'd39; 
32'd1220: dataIn1 = 32'd25; 
32'd1221: dataIn1 = 32'd8; 
32'd1222: dataIn1 = 32'd13; 
32'd1223: dataIn1 = 32'd23; 
32'd1224: dataIn1 = 32'd53; 
32'd1225: dataIn1 = 32'd62; 
32'd1226: dataIn1 = 32'd26; 
32'd1227: dataIn1 = 32'd0; 
32'd1228: dataIn1 = 32'd57; 
32'd1229: dataIn1 = 32'd15; 
32'd1230: dataIn1 = 32'd3; 
32'd1231: dataIn1 = 32'd51; 
32'd1232: dataIn1 = 32'd14; 
32'd1233: dataIn1 = 32'd1; 
32'd1234: dataIn1 = 32'd1; 
32'd1235: dataIn1 = 32'd38; 
32'd1236: dataIn1 = 32'd26; 
32'd1237: dataIn1 = 32'd57; 
32'd1238: dataIn1 = 32'd50; 
32'd1239: dataIn1 = 32'd47; 
32'd1240: dataIn1 = 32'd36; 
32'd1241: dataIn1 = 32'd44; 
32'd1242: dataIn1 = 32'd10; 
32'd1243: dataIn1 = 32'd50; 
32'd1244: dataIn1 = 32'd49; 
32'd1245: dataIn1 = 32'd1; 
32'd1246: dataIn1 = 32'd31; 
32'd1247: dataIn1 = 32'd22; 
32'd1248: dataIn1 = 32'd41; 
32'd1249: dataIn1 = 32'd46; 
32'd1250: dataIn1 = 32'd21; 
32'd1251: dataIn1 = 32'd58; 
32'd1252: dataIn1 = 32'd37; 
32'd1253: dataIn1 = 32'd37; 
32'd1254: dataIn1 = 32'd59; 
32'd1255: dataIn1 = 32'd8; 
32'd1256: dataIn1 = 32'd19; 
32'd1257: dataIn1 = 32'd60; 
32'd1258: dataIn1 = 32'd41; 
32'd1259: dataIn1 = 32'd32; 
32'd1260: dataIn1 = 32'd16; 
32'd1261: dataIn1 = 32'd20; 
32'd1262: dataIn1 = 32'd45; 
32'd1263: dataIn1 = 32'd54; 
32'd1264: dataIn1 = 32'd2; 
32'd1265: dataIn1 = 32'd43; 
32'd1266: dataIn1 = 32'd16; 
32'd1267: dataIn1 = 32'd38; 
32'd1268: dataIn1 = 32'd27; 
32'd1269: dataIn1 = 32'd62; 
32'd1270: dataIn1 = 32'd51; 
32'd1271: dataIn1 = 32'd17; 
32'd1272: dataIn1 = 32'd2; 
32'd1273: dataIn1 = 32'd6; 
32'd1274: dataIn1 = 32'd40; 
32'd1275: dataIn1 = 32'd61; 
32'd1276: dataIn1 = 32'd20; 
32'd1277: dataIn1 = 32'd49; 
32'd1278: dataIn1 = 32'd30; 
32'd1279: dataIn1 = 32'd17; 
32'd1280: dataIn1 = 32'd33; 
32'd1281: dataIn1 = 32'd35; 
32'd1282: dataIn1 = 32'd37; 
32'd1283: dataIn1 = 32'd58; 
32'd1284: dataIn1 = 32'd4; 
32'd1285: dataIn1 = 32'd7; 
32'd1286: dataIn1 = 32'd44; 
32'd1287: dataIn1 = 32'd20; 
32'd1288: dataIn1 = 32'd16; 
32'd1289: dataIn1 = 32'd55; 
32'd1290: dataIn1 = 32'd36; 
32'd1291: dataIn1 = 32'd3; 
32'd1292: dataIn1 = 32'd6; 
32'd1293: dataIn1 = 32'd45; 
32'd1294: dataIn1 = 32'd47; 
32'd1295: dataIn1 = 32'd47; 
32'd1296: dataIn1 = 32'd13; 
32'd1297: dataIn1 = 32'd36; 
32'd1298: dataIn1 = 32'd53; 
32'd1299: dataIn1 = 32'd26; 
32'd1300: dataIn1 = 32'd42; 
32'd1301: dataIn1 = 32'd18; 
32'd1302: dataIn1 = 32'd61; 
32'd1303: dataIn1 = 32'd32; 
32'd1304: dataIn1 = 32'd54; 
32'd1305: dataIn1 = 32'd61; 
32'd1306: dataIn1 = 32'd4; 
32'd1307: dataIn1 = 32'd22; 
32'd1308: dataIn1 = 32'd44; 
32'd1309: dataIn1 = 32'd7; 
32'd1310: dataIn1 = 32'd42; 
32'd1311: dataIn1 = 32'd63; 
32'd1312: dataIn1 = 32'd7; 
32'd1313: dataIn1 = 32'd18; 
32'd1314: dataIn1 = 32'd52; 
32'd1315: dataIn1 = 32'd35; 
32'd1316: dataIn1 = 32'd55; 
32'd1317: dataIn1 = 32'd0; 
32'd1318: dataIn1 = 32'd34; 
32'd1319: dataIn1 = 32'd47; 
32'd1320: dataIn1 = 32'd6; 
32'd1321: dataIn1 = 32'd36; 
32'd1322: dataIn1 = 32'd18; 
32'd1323: dataIn1 = 32'd18; 
32'd1324: dataIn1 = 32'd38; 
32'd1325: dataIn1 = 32'd34; 
32'd1326: dataIn1 = 32'd59; 
32'd1327: dataIn1 = 32'd55; 
32'd1328: dataIn1 = 32'd47; 
32'd1329: dataIn1 = 32'd58; 
32'd1330: dataIn1 = 32'd20; 
32'd1331: dataIn1 = 32'd15; 
32'd1332: dataIn1 = 32'd52; 
32'd1333: dataIn1 = 32'd48; 
32'd1334: dataIn1 = 32'd48; 
32'd1335: dataIn1 = 32'd60; 
32'd1336: dataIn1 = 32'd31; 
32'd1337: dataIn1 = 32'd27; 
32'd1338: dataIn1 = 32'd9; 
32'd1339: dataIn1 = 32'd39; 
32'd1340: dataIn1 = 32'd40; 
32'd1341: dataIn1 = 32'd4; 
32'd1342: dataIn1 = 32'd58; 
32'd1343: dataIn1 = 32'd5; 
32'd1344: dataIn1 = 32'd27; 
32'd1345: dataIn1 = 32'd3; 
32'd1346: dataIn1 = 32'd37; 
32'd1347: dataIn1 = 32'd38; 
32'd1348: dataIn1 = 32'd48; 
32'd1349: dataIn1 = 32'd13; 
32'd1350: dataIn1 = 32'd35; 
32'd1351: dataIn1 = 32'd3; 
32'd1352: dataIn1 = 32'd14; 
32'd1353: dataIn1 = 32'd46; 
32'd1354: dataIn1 = 32'd63; 
32'd1355: dataIn1 = 32'd40; 
32'd1356: dataIn1 = 32'd57; 
32'd1357: dataIn1 = 32'd62; 
32'd1358: dataIn1 = 32'd32; 
32'd1359: dataIn1 = 32'd50; 
32'd1360: dataIn1 = 32'd42; 
32'd1361: dataIn1 = 32'd18; 
32'd1362: dataIn1 = 32'd61; 
32'd1363: dataIn1 = 32'd37; 
32'd1364: dataIn1 = 32'd23; 
32'd1365: dataIn1 = 32'd57; 
32'd1366: dataIn1 = 32'd42; 
32'd1367: dataIn1 = 32'd4; 
32'd1368: dataIn1 = 32'd33; 
32'd1369: dataIn1 = 32'd50; 
32'd1370: dataIn1 = 32'd2; 
32'd1371: dataIn1 = 32'd14; 
32'd1372: dataIn1 = 32'd55; 
32'd1373: dataIn1 = 32'd54; 
32'd1374: dataIn1 = 32'd26; 
32'd1375: dataIn1 = 32'd31; 
32'd1376: dataIn1 = 32'd17; 
32'd1377: dataIn1 = 32'd9; 
32'd1378: dataIn1 = 32'd28; 
32'd1379: dataIn1 = 32'd51; 
32'd1380: dataIn1 = 32'd18; 
32'd1381: dataIn1 = 32'd48; 
32'd1382: dataIn1 = 32'd18; 
32'd1383: dataIn1 = 32'd6; 
32'd1384: dataIn1 = 32'd19; 
32'd1385: dataIn1 = 32'd16; 
32'd1386: dataIn1 = 32'd21; 
32'd1387: dataIn1 = 32'd42; 
32'd1388: dataIn1 = 32'd1; 
32'd1389: dataIn1 = 32'd17; 
32'd1390: dataIn1 = 32'd18; 
32'd1391: dataIn1 = 32'd26; 
32'd1392: dataIn1 = 32'd18; 
32'd1393: dataIn1 = 32'd25; 
32'd1394: dataIn1 = 32'd0; 
32'd1395: dataIn1 = 32'd60; 
32'd1396: dataIn1 = 32'd1; 
32'd1397: dataIn1 = 32'd51; 
32'd1398: dataIn1 = 32'd21; 
32'd1399: dataIn1 = 32'd14; 
32'd1400: dataIn1 = 32'd63; 
32'd1401: dataIn1 = 32'd44; 
32'd1402: dataIn1 = 32'd16; 
32'd1403: dataIn1 = 32'd10; 
32'd1404: dataIn1 = 32'd33; 
32'd1405: dataIn1 = 32'd59; 
32'd1406: dataIn1 = 32'd17; 
32'd1407: dataIn1 = 32'd35; 
32'd1408: dataIn1 = 32'd7; 
32'd1409: dataIn1 = 32'd48; 
32'd1410: dataIn1 = 32'd58; 
32'd1411: dataIn1 = 32'd32; 
32'd1412: dataIn1 = 32'd28; 
32'd1413: dataIn1 = 32'd52; 
32'd1414: dataIn1 = 32'd30; 
32'd1415: dataIn1 = 32'd53; 
32'd1416: dataIn1 = 32'd23; 
32'd1417: dataIn1 = 32'd32; 
32'd1418: dataIn1 = 32'd44; 
32'd1419: dataIn1 = 32'd48; 
32'd1420: dataIn1 = 32'd19; 
32'd1421: dataIn1 = 32'd9; 
32'd1422: dataIn1 = 32'd33; 
32'd1423: dataIn1 = 32'd8; 
32'd1424: dataIn1 = 32'd37; 
32'd1425: dataIn1 = 32'd27; 
32'd1426: dataIn1 = 32'd12; 
32'd1427: dataIn1 = 32'd0; 
32'd1428: dataIn1 = 32'd21; 
32'd1429: dataIn1 = 32'd51; 
32'd1430: dataIn1 = 32'd15; 
32'd1431: dataIn1 = 32'd51; 
32'd1432: dataIn1 = 32'd1; 
32'd1433: dataIn1 = 32'd52; 
32'd1434: dataIn1 = 32'd31; 
32'd1435: dataIn1 = 32'd15; 
32'd1436: dataIn1 = 32'd9; 
32'd1437: dataIn1 = 32'd12; 
32'd1438: dataIn1 = 32'd62; 
32'd1439: dataIn1 = 32'd9; 
32'd1440: dataIn1 = 32'd29; 
32'd1441: dataIn1 = 32'd29; 
32'd1442: dataIn1 = 32'd54; 
32'd1443: dataIn1 = 32'd43; 
32'd1444: dataIn1 = 32'd59; 
32'd1445: dataIn1 = 32'd2; 
32'd1446: dataIn1 = 32'd26; 
32'd1447: dataIn1 = 32'd50; 
32'd1448: dataIn1 = 32'd27; 
32'd1449: dataIn1 = 32'd6; 
32'd1450: dataIn1 = 32'd39; 
32'd1451: dataIn1 = 32'd12; 
32'd1452: dataIn1 = 32'd41; 
32'd1453: dataIn1 = 32'd22; 
32'd1454: dataIn1 = 32'd33; 
32'd1455: dataIn1 = 32'd32; 
32'd1456: dataIn1 = 32'd39; 
32'd1457: dataIn1 = 32'd21; 
32'd1458: dataIn1 = 32'd53; 
32'd1459: dataIn1 = 32'd47; 
32'd1460: dataIn1 = 32'd21; 
32'd1461: dataIn1 = 32'd1; 
32'd1462: dataIn1 = 32'd29; 
32'd1463: dataIn1 = 32'd38; 
32'd1464: dataIn1 = 32'd29; 
32'd1465: dataIn1 = 32'd50; 
32'd1466: dataIn1 = 32'd59; 
32'd1467: dataIn1 = 32'd8; 
32'd1468: dataIn1 = 32'd36; 
32'd1469: dataIn1 = 32'd57; 
32'd1470: dataIn1 = 32'd6; 
32'd1471: dataIn1 = 32'd61; 
32'd1472: dataIn1 = 32'd12; 
32'd1473: dataIn1 = 32'd3; 
32'd1474: dataIn1 = 32'd28; 
32'd1475: dataIn1 = 32'd17; 
32'd1476: dataIn1 = 32'd42; 
32'd1477: dataIn1 = 32'd7; 
32'd1478: dataIn1 = 32'd48; 
32'd1479: dataIn1 = 32'd51; 
32'd1480: dataIn1 = 32'd13; 
32'd1481: dataIn1 = 32'd51; 
32'd1482: dataIn1 = 32'd60; 
32'd1483: dataIn1 = 32'd6; 
32'd1484: dataIn1 = 32'd3; 
32'd1485: dataIn1 = 32'd15; 
32'd1486: dataIn1 = 32'd61; 
32'd1487: dataIn1 = 32'd5; 
32'd1488: dataIn1 = 32'd23; 
32'd1489: dataIn1 = 32'd20; 
32'd1490: dataIn1 = 32'd18; 
32'd1491: dataIn1 = 32'd51; 
32'd1492: dataIn1 = 32'd47; 
32'd1493: dataIn1 = 32'd57; 
32'd1494: dataIn1 = 32'd13; 
32'd1495: dataIn1 = 32'd56; 
32'd1496: dataIn1 = 32'd37; 
32'd1497: dataIn1 = 32'd39; 
32'd1498: dataIn1 = 32'd27; 
32'd1499: dataIn1 = 32'd37; 
32'd1500: dataIn1 = 32'd33; 
32'd1501: dataIn1 = 32'd55; 
32'd1502: dataIn1 = 32'd36; 
32'd1503: dataIn1 = 32'd61; 
32'd1504: dataIn1 = 32'd28; 
32'd1505: dataIn1 = 32'd47; 
32'd1506: dataIn1 = 32'd11; 
32'd1507: dataIn1 = 32'd47; 
32'd1508: dataIn1 = 32'd1; 
32'd1509: dataIn1 = 32'd25; 
32'd1510: dataIn1 = 32'd32; 
32'd1511: dataIn1 = 32'd43; 
32'd1512: dataIn1 = 32'd15; 
32'd1513: dataIn1 = 32'd37; 
32'd1514: dataIn1 = 32'd60; 
32'd1515: dataIn1 = 32'd14; 
32'd1516: dataIn1 = 32'd54; 
32'd1517: dataIn1 = 32'd25; 
32'd1518: dataIn1 = 32'd20; 
32'd1519: dataIn1 = 32'd2; 
32'd1520: dataIn1 = 32'd1; 
32'd1521: dataIn1 = 32'd58; 
32'd1522: dataIn1 = 32'd48; 
32'd1523: dataIn1 = 32'd3; 
32'd1524: dataIn1 = 32'd54; 
32'd1525: dataIn1 = 32'd36; 
32'd1526: dataIn1 = 32'd28; 
32'd1527: dataIn1 = 32'd57; 
32'd1528: dataIn1 = 32'd5; 
32'd1529: dataIn1 = 32'd19; 
32'd1530: dataIn1 = 32'd50; 
32'd1531: dataIn1 = 32'd33; 
32'd1532: dataIn1 = 32'd47; 
32'd1533: dataIn1 = 32'd17; 
32'd1534: dataIn1 = 32'd54; 
32'd1535: dataIn1 = 32'd4; 
32'd1536: dataIn1 = 32'd26; 
32'd1537: dataIn1 = 32'd37; 
32'd1538: dataIn1 = 32'd58; 
32'd1539: dataIn1 = 32'd59; 
32'd1540: dataIn1 = 32'd16; 
32'd1541: dataIn1 = 32'd9; 
32'd1542: dataIn1 = 32'd55; 
32'd1543: dataIn1 = 32'd10; 
32'd1544: dataIn1 = 32'd22; 
32'd1545: dataIn1 = 32'd38; 
32'd1546: dataIn1 = 32'd38; 
32'd1547: dataIn1 = 32'd58; 
32'd1548: dataIn1 = 32'd56; 
32'd1549: dataIn1 = 32'd21; 
32'd1550: dataIn1 = 32'd0; 
32'd1551: dataIn1 = 32'd23; 
32'd1552: dataIn1 = 32'd52; 
32'd1553: dataIn1 = 32'd1; 
32'd1554: dataIn1 = 32'd56; 
32'd1555: dataIn1 = 32'd32; 
32'd1556: dataIn1 = 32'd1; 
32'd1557: dataIn1 = 32'd58; 
32'd1558: dataIn1 = 32'd35; 
32'd1559: dataIn1 = 32'd49; 
32'd1560: dataIn1 = 32'd9; 
32'd1561: dataIn1 = 32'd54; 
32'd1562: dataIn1 = 32'd7; 
32'd1563: dataIn1 = 32'd46; 
32'd1564: dataIn1 = 32'd39; 
32'd1565: dataIn1 = 32'd28; 
32'd1566: dataIn1 = 32'd3; 
32'd1567: dataIn1 = 32'd54; 
32'd1568: dataIn1 = 32'd44; 
32'd1569: dataIn1 = 32'd0; 
32'd1570: dataIn1 = 32'd13; 
32'd1571: dataIn1 = 32'd54; 
32'd1572: dataIn1 = 32'd52; 
32'd1573: dataIn1 = 32'd57; 
32'd1574: dataIn1 = 32'd11; 
32'd1575: dataIn1 = 32'd5; 
32'd1576: dataIn1 = 32'd46; 
32'd1577: dataIn1 = 32'd39; 
32'd1578: dataIn1 = 32'd32; 
32'd1579: dataIn1 = 32'd29; 
32'd1580: dataIn1 = 32'd14; 
32'd1581: dataIn1 = 32'd43; 
32'd1582: dataIn1 = 32'd14; 
32'd1583: dataIn1 = 32'd10; 
32'd1584: dataIn1 = 32'd24; 
32'd1585: dataIn1 = 32'd40; 
32'd1586: dataIn1 = 32'd57; 
32'd1587: dataIn1 = 32'd46; 
32'd1588: dataIn1 = 32'd4; 
32'd1589: dataIn1 = 32'd29; 
32'd1590: dataIn1 = 32'd45; 
32'd1591: dataIn1 = 32'd32; 
32'd1592: dataIn1 = 32'd40; 
32'd1593: dataIn1 = 32'd45; 
32'd1594: dataIn1 = 32'd44; 
32'd1595: dataIn1 = 32'd33; 
32'd1596: dataIn1 = 32'd53; 
32'd1597: dataIn1 = 32'd29; 
32'd1598: dataIn1 = 32'd40; 
32'd1599: dataIn1 = 32'd50; 
32'd1600: dataIn1 = 32'd2; 
32'd1601: dataIn1 = 32'd10; 
32'd1602: dataIn1 = 32'd56; 
32'd1603: dataIn1 = 32'd63; 
32'd1604: dataIn1 = 32'd36; 
32'd1605: dataIn1 = 32'd22; 
32'd1606: dataIn1 = 32'd23; 
32'd1607: dataIn1 = 32'd12; 
32'd1608: dataIn1 = 32'd16; 
32'd1609: dataIn1 = 32'd8; 
32'd1610: dataIn1 = 32'd4; 
32'd1611: dataIn1 = 32'd4; 
32'd1612: dataIn1 = 32'd29; 
32'd1613: dataIn1 = 32'd38; 
32'd1614: dataIn1 = 32'd52; 
32'd1615: dataIn1 = 32'd28; 
32'd1616: dataIn1 = 32'd29; 
32'd1617: dataIn1 = 32'd24; 
32'd1618: dataIn1 = 32'd60; 
32'd1619: dataIn1 = 32'd33; 
32'd1620: dataIn1 = 32'd11; 
32'd1621: dataIn1 = 32'd42; 
32'd1622: dataIn1 = 32'd4; 
32'd1623: dataIn1 = 32'd47; 
32'd1624: dataIn1 = 32'd20; 
32'd1625: dataIn1 = 32'd46; 
32'd1626: dataIn1 = 32'd32; 
32'd1627: dataIn1 = 32'd39; 
32'd1628: dataIn1 = 32'd15; 
32'd1629: dataIn1 = 32'd30; 
32'd1630: dataIn1 = 32'd24; 
32'd1631: dataIn1 = 32'd0; 
32'd1632: dataIn1 = 32'd30; 
32'd1633: dataIn1 = 32'd43; 
32'd1634: dataIn1 = 32'd17; 
32'd1635: dataIn1 = 32'd47; 
32'd1636: dataIn1 = 32'd55; 
32'd1637: dataIn1 = 32'd61; 
32'd1638: dataIn1 = 32'd15; 
32'd1639: dataIn1 = 32'd9; 
32'd1640: dataIn1 = 32'd14; 
32'd1641: dataIn1 = 32'd58; 
32'd1642: dataIn1 = 32'd37; 
32'd1643: dataIn1 = 32'd59; 
32'd1644: dataIn1 = 32'd38; 
32'd1645: dataIn1 = 32'd10; 
32'd1646: dataIn1 = 32'd12; 
32'd1647: dataIn1 = 32'd21; 
32'd1648: dataIn1 = 32'd13; 
32'd1649: dataIn1 = 32'd42; 
32'd1650: dataIn1 = 32'd43; 
32'd1651: dataIn1 = 32'd62; 
32'd1652: dataIn1 = 32'd13; 
32'd1653: dataIn1 = 32'd56; 
32'd1654: dataIn1 = 32'd25; 
32'd1655: dataIn1 = 32'd6; 
32'd1656: dataIn1 = 32'd54; 
32'd1657: dataIn1 = 32'd25; 
32'd1658: dataIn1 = 32'd10; 
32'd1659: dataIn1 = 32'd63; 
32'd1660: dataIn1 = 32'd27; 
32'd1661: dataIn1 = 32'd38; 
32'd1662: dataIn1 = 32'd57; 
32'd1663: dataIn1 = 32'd37; 
32'd1664: dataIn1 = 32'd5; 
32'd1665: dataIn1 = 32'd5; 
32'd1666: dataIn1 = 32'd10; 
32'd1667: dataIn1 = 32'd28; 
32'd1668: dataIn1 = 32'd34; 
32'd1669: dataIn1 = 32'd46; 
32'd1670: dataIn1 = 32'd17; 
32'd1671: dataIn1 = 32'd14; 
32'd1672: dataIn1 = 32'd24; 
32'd1673: dataIn1 = 32'd7; 
32'd1674: dataIn1 = 32'd57; 
32'd1675: dataIn1 = 32'd5; 
32'd1676: dataIn1 = 32'd51; 
32'd1677: dataIn1 = 32'd21; 
32'd1678: dataIn1 = 32'd16; 
32'd1679: dataIn1 = 32'd51; 
32'd1680: dataIn1 = 32'd1; 
32'd1681: dataIn1 = 32'd25; 
32'd1682: dataIn1 = 32'd14; 
32'd1683: dataIn1 = 32'd37; 
32'd1684: dataIn1 = 32'd8; 
32'd1685: dataIn1 = 32'd2; 
32'd1686: dataIn1 = 32'd43; 
32'd1687: dataIn1 = 32'd0; 
32'd1688: dataIn1 = 32'd20; 
32'd1689: dataIn1 = 32'd46; 
32'd1690: dataIn1 = 32'd21; 
32'd1691: dataIn1 = 32'd59; 
32'd1692: dataIn1 = 32'd63; 
32'd1693: dataIn1 = 32'd40; 
32'd1694: dataIn1 = 32'd34; 
32'd1695: dataIn1 = 32'd35; 
32'd1696: dataIn1 = 32'd6; 
32'd1697: dataIn1 = 32'd24; 
32'd1698: dataIn1 = 32'd40; 
32'd1699: dataIn1 = 32'd8; 
32'd1700: dataIn1 = 32'd17; 
32'd1701: dataIn1 = 32'd24; 
32'd1702: dataIn1 = 32'd38; 
32'd1703: dataIn1 = 32'd49; 
32'd1704: dataIn1 = 32'd39; 
32'd1705: dataIn1 = 32'd35; 
32'd1706: dataIn1 = 32'd21; 
32'd1707: dataIn1 = 32'd6; 
32'd1708: dataIn1 = 32'd43; 
32'd1709: dataIn1 = 32'd47; 
32'd1710: dataIn1 = 32'd38; 
32'd1711: dataIn1 = 32'd52; 
32'd1712: dataIn1 = 32'd6; 
32'd1713: dataIn1 = 32'd6; 
32'd1714: dataIn1 = 32'd16; 
32'd1715: dataIn1 = 32'd4; 
32'd1716: dataIn1 = 32'd50; 
32'd1717: dataIn1 = 32'd39; 
32'd1718: dataIn1 = 32'd19; 
32'd1719: dataIn1 = 32'd39; 
32'd1720: dataIn1 = 32'd48; 
32'd1721: dataIn1 = 32'd0; 
32'd1722: dataIn1 = 32'd56; 
32'd1723: dataIn1 = 32'd4; 
32'd1724: dataIn1 = 32'd20; 
32'd1725: dataIn1 = 32'd13; 
32'd1726: dataIn1 = 32'd4; 
32'd1727: dataIn1 = 32'd20; 
32'd1728: dataIn1 = 32'd35; 
32'd1729: dataIn1 = 32'd62; 
32'd1730: dataIn1 = 32'd26; 
32'd1731: dataIn1 = 32'd12; 
32'd1732: dataIn1 = 32'd13; 
32'd1733: dataIn1 = 32'd28; 
32'd1734: dataIn1 = 32'd33; 
32'd1735: dataIn1 = 32'd31; 
32'd1736: dataIn1 = 32'd35; 
32'd1737: dataIn1 = 32'd17; 
32'd1738: dataIn1 = 32'd52; 
32'd1739: dataIn1 = 32'd10; 
32'd1740: dataIn1 = 32'd21; 
32'd1741: dataIn1 = 32'd1; 
32'd1742: dataIn1 = 32'd25; 
32'd1743: dataIn1 = 32'd3; 
32'd1744: dataIn1 = 32'd6; 
32'd1745: dataIn1 = 32'd15; 
32'd1746: dataIn1 = 32'd8; 
32'd1747: dataIn1 = 32'd16; 
32'd1748: dataIn1 = 32'd4; 
32'd1749: dataIn1 = 32'd53; 
32'd1750: dataIn1 = 32'd16; 
32'd1751: dataIn1 = 32'd61; 
32'd1752: dataIn1 = 32'd27; 
32'd1753: dataIn1 = 32'd13; 
32'd1754: dataIn1 = 32'd21; 
32'd1755: dataIn1 = 32'd29; 
32'd1756: dataIn1 = 32'd4; 
32'd1757: dataIn1 = 32'd55; 
32'd1758: dataIn1 = 32'd35; 
32'd1759: dataIn1 = 32'd0; 
32'd1760: dataIn1 = 32'd1; 
32'd1761: dataIn1 = 32'd51; 
32'd1762: dataIn1 = 32'd34; 
32'd1763: dataIn1 = 32'd9; 
32'd1764: dataIn1 = 32'd45; 
32'd1765: dataIn1 = 32'd63; 
32'd1766: dataIn1 = 32'd23; 
32'd1767: dataIn1 = 32'd56; 
32'd1768: dataIn1 = 32'd21; 
32'd1769: dataIn1 = 32'd34; 
32'd1770: dataIn1 = 32'd12; 
32'd1771: dataIn1 = 32'd1; 
32'd1772: dataIn1 = 32'd48; 
32'd1773: dataIn1 = 32'd28; 
32'd1774: dataIn1 = 32'd22; 
32'd1775: dataIn1 = 32'd31; 
32'd1776: dataIn1 = 32'd55; 
32'd1777: dataIn1 = 32'd56; 
32'd1778: dataIn1 = 32'd34; 
32'd1779: dataIn1 = 32'd24; 
32'd1780: dataIn1 = 32'd49; 
32'd1781: dataIn1 = 32'd61; 
32'd1782: dataIn1 = 32'd58; 
32'd1783: dataIn1 = 32'd21; 
32'd1784: dataIn1 = 32'd62; 
32'd1785: dataIn1 = 32'd56; 
32'd1786: dataIn1 = 32'd45; 
32'd1787: dataIn1 = 32'd4; 
32'd1788: dataIn1 = 32'd24; 
32'd1789: dataIn1 = 32'd4; 
32'd1790: dataIn1 = 32'd10; 
32'd1791: dataIn1 = 32'd57; 
32'd1792: dataIn1 = 32'd19; 
32'd1793: dataIn1 = 32'd51; 
32'd1794: dataIn1 = 32'd19; 
32'd1795: dataIn1 = 32'd59; 
32'd1796: dataIn1 = 32'd40; 
32'd1797: dataIn1 = 32'd42; 
32'd1798: dataIn1 = 32'd2; 
32'd1799: dataIn1 = 32'd49; 
32'd1800: dataIn1 = 32'd38; 
32'd1801: dataIn1 = 32'd0; 
32'd1802: dataIn1 = 32'd33; 
32'd1803: dataIn1 = 32'd59; 
32'd1804: dataIn1 = 32'd19; 
32'd1805: dataIn1 = 32'd53; 
32'd1806: dataIn1 = 32'd15; 
32'd1807: dataIn1 = 32'd25; 
32'd1808: dataIn1 = 32'd12; 
32'd1809: dataIn1 = 32'd54; 
32'd1810: dataIn1 = 32'd31; 
32'd1811: dataIn1 = 32'd27; 
32'd1812: dataIn1 = 32'd45; 
32'd1813: dataIn1 = 32'd52; 
32'd1814: dataIn1 = 32'd45; 
32'd1815: dataIn1 = 32'd49; 
32'd1816: dataIn1 = 32'd61; 
32'd1817: dataIn1 = 32'd22; 
32'd1818: dataIn1 = 32'd12; 
32'd1819: dataIn1 = 32'd41; 
32'd1820: dataIn1 = 32'd53; 
32'd1821: dataIn1 = 32'd54; 
32'd1822: dataIn1 = 32'd36; 
32'd1823: dataIn1 = 32'd11; 
32'd1824: dataIn1 = 32'd53; 
32'd1825: dataIn1 = 32'd61; 
32'd1826: dataIn1 = 32'd12; 
32'd1827: dataIn1 = 32'd46; 
32'd1828: dataIn1 = 32'd17; 
32'd1829: dataIn1 = 32'd51; 
32'd1830: dataIn1 = 32'd25; 
32'd1831: dataIn1 = 32'd2; 
32'd1832: dataIn1 = 32'd13; 
32'd1833: dataIn1 = 32'd25; 
32'd1834: dataIn1 = 32'd36; 
32'd1835: dataIn1 = 32'd51; 
32'd1836: dataIn1 = 32'd50; 
32'd1837: dataIn1 = 32'd15; 
32'd1838: dataIn1 = 32'd3; 
32'd1839: dataIn1 = 32'd25; 
32'd1840: dataIn1 = 32'd40; 
32'd1841: dataIn1 = 32'd41; 
32'd1842: dataIn1 = 32'd56; 
32'd1843: dataIn1 = 32'd4; 
32'd1844: dataIn1 = 32'd53; 
32'd1845: dataIn1 = 32'd5; 
32'd1846: dataIn1 = 32'd41; 
32'd1847: dataIn1 = 32'd51; 
32'd1848: dataIn1 = 32'd47; 
32'd1849: dataIn1 = 32'd40; 
32'd1850: dataIn1 = 32'd38; 
32'd1851: dataIn1 = 32'd57; 
32'd1852: dataIn1 = 32'd25; 
32'd1853: dataIn1 = 32'd30; 
32'd1854: dataIn1 = 32'd6; 
32'd1855: dataIn1 = 32'd13; 
32'd1856: dataIn1 = 32'd24; 
32'd1857: dataIn1 = 32'd41; 
32'd1858: dataIn1 = 32'd42; 
32'd1859: dataIn1 = 32'd28; 
32'd1860: dataIn1 = 32'd41; 
32'd1861: dataIn1 = 32'd23; 
32'd1862: dataIn1 = 32'd56; 
32'd1863: dataIn1 = 32'd35; 
32'd1864: dataIn1 = 32'd39; 
32'd1865: dataIn1 = 32'd47; 
32'd1866: dataIn1 = 32'd31; 
32'd1867: dataIn1 = 32'd17; 
32'd1868: dataIn1 = 32'd32; 
32'd1869: dataIn1 = 32'd54; 
32'd1870: dataIn1 = 32'd13; 
32'd1871: dataIn1 = 32'd58; 
32'd1872: dataIn1 = 32'd40; 
32'd1873: dataIn1 = 32'd1; 
32'd1874: dataIn1 = 32'd14; 
32'd1875: dataIn1 = 32'd63; 
32'd1876: dataIn1 = 32'd45; 
32'd1877: dataIn1 = 32'd29; 
32'd1878: dataIn1 = 32'd26; 
32'd1879: dataIn1 = 32'd40; 
32'd1880: dataIn1 = 32'd30; 
32'd1881: dataIn1 = 32'd36; 
32'd1882: dataIn1 = 32'd12; 
32'd1883: dataIn1 = 32'd59; 
32'd1884: dataIn1 = 32'd29; 
32'd1885: dataIn1 = 32'd51; 
32'd1886: dataIn1 = 32'd48; 
32'd1887: dataIn1 = 32'd27; 
32'd1888: dataIn1 = 32'd54; 
32'd1889: dataIn1 = 32'd5; 
32'd1890: dataIn1 = 32'd6; 
32'd1891: dataIn1 = 32'd62; 
32'd1892: dataIn1 = 32'd41; 
32'd1893: dataIn1 = 32'd55; 
32'd1894: dataIn1 = 32'd23; 
32'd1895: dataIn1 = 32'd11; 
32'd1896: dataIn1 = 32'd39; 
32'd1897: dataIn1 = 32'd25; 
32'd1898: dataIn1 = 32'd24; 
32'd1899: dataIn1 = 32'd8; 
32'd1900: dataIn1 = 32'd3; 
32'd1901: dataIn1 = 32'd51; 
32'd1902: dataIn1 = 32'd62; 
32'd1903: dataIn1 = 32'd4; 
32'd1904: dataIn1 = 32'd22; 
32'd1905: dataIn1 = 32'd63; 
32'd1906: dataIn1 = 32'd21; 
32'd1907: dataIn1 = 32'd0; 
32'd1908: dataIn1 = 32'd9; 
32'd1909: dataIn1 = 32'd59; 
32'd1910: dataIn1 = 32'd37; 
32'd1911: dataIn1 = 32'd47; 
32'd1912: dataIn1 = 32'd26; 
32'd1913: dataIn1 = 32'd23; 
32'd1914: dataIn1 = 32'd11; 
32'd1915: dataIn1 = 32'd56; 
32'd1916: dataIn1 = 32'd57; 
32'd1917: dataIn1 = 32'd53; 
32'd1918: dataIn1 = 32'd59; 
32'd1919: dataIn1 = 32'd48; 
32'd1920: dataIn1 = 32'd50; 
32'd1921: dataIn1 = 32'd19; 
32'd1922: dataIn1 = 32'd1; 
32'd1923: dataIn1 = 32'd50; 
32'd1924: dataIn1 = 32'd38; 
32'd1925: dataIn1 = 32'd4; 
32'd1926: dataIn1 = 32'd44; 
32'd1927: dataIn1 = 32'd13; 
32'd1928: dataIn1 = 32'd63; 
32'd1929: dataIn1 = 32'd4; 
32'd1930: dataIn1 = 32'd20; 
32'd1931: dataIn1 = 32'd58; 
32'd1932: dataIn1 = 32'd6; 
32'd1933: dataIn1 = 32'd11; 
32'd1934: dataIn1 = 32'd62; 
32'd1935: dataIn1 = 32'd26; 
32'd1936: dataIn1 = 32'd28; 
32'd1937: dataIn1 = 32'd53; 
32'd1938: dataIn1 = 32'd15; 
32'd1939: dataIn1 = 32'd35; 
32'd1940: dataIn1 = 32'd1; 
32'd1941: dataIn1 = 32'd9; 
32'd1942: dataIn1 = 32'd22; 
32'd1943: dataIn1 = 32'd4; 
32'd1944: dataIn1 = 32'd10; 
32'd1945: dataIn1 = 32'd9; 
32'd1946: dataIn1 = 32'd28; 
32'd1947: dataIn1 = 32'd52; 
32'd1948: dataIn1 = 32'd30; 
32'd1949: dataIn1 = 32'd12; 
32'd1950: dataIn1 = 32'd28; 
32'd1951: dataIn1 = 32'd54; 
32'd1952: dataIn1 = 32'd44; 
32'd1953: dataIn1 = 32'd12; 
32'd1954: dataIn1 = 32'd36; 
32'd1955: dataIn1 = 32'd16; 
32'd1956: dataIn1 = 32'd30; 
32'd1957: dataIn1 = 32'd46; 
32'd1958: dataIn1 = 32'd11; 
32'd1959: dataIn1 = 32'd55; 
32'd1960: dataIn1 = 32'd11; 
32'd1961: dataIn1 = 32'd28; 
32'd1962: dataIn1 = 32'd58; 
32'd1963: dataIn1 = 32'd27; 
32'd1964: dataIn1 = 32'd57; 
32'd1965: dataIn1 = 32'd32; 
32'd1966: dataIn1 = 32'd42; 
32'd1967: dataIn1 = 32'd54; 
32'd1968: dataIn1 = 32'd7; 
32'd1969: dataIn1 = 32'd23; 
32'd1970: dataIn1 = 32'd1; 
32'd1971: dataIn1 = 32'd4; 
32'd1972: dataIn1 = 32'd53; 
32'd1973: dataIn1 = 32'd30; 
32'd1974: dataIn1 = 32'd37; 
32'd1975: dataIn1 = 32'd51; 
32'd1976: dataIn1 = 32'd19; 
32'd1977: dataIn1 = 32'd63; 
32'd1978: dataIn1 = 32'd19; 
32'd1979: dataIn1 = 32'd59; 
32'd1980: dataIn1 = 32'd47; 
32'd1981: dataIn1 = 32'd16; 
32'd1982: dataIn1 = 32'd12; 
32'd1983: dataIn1 = 32'd55; 
32'd1984: dataIn1 = 32'd36; 
32'd1985: dataIn1 = 32'd4; 
32'd1986: dataIn1 = 32'd3; 
32'd1987: dataIn1 = 32'd10; 
32'd1988: dataIn1 = 32'd14; 
32'd1989: dataIn1 = 32'd51; 
32'd1990: dataIn1 = 32'd28; 
32'd1991: dataIn1 = 32'd14; 
32'd1992: dataIn1 = 32'd28; 
32'd1993: dataIn1 = 32'd38; 
32'd1994: dataIn1 = 32'd46; 
32'd1995: dataIn1 = 32'd5; 
32'd1996: dataIn1 = 32'd56; 
32'd1997: dataIn1 = 32'd42; 
32'd1998: dataIn1 = 32'd51; 
32'd1999: dataIn1 = 32'd15; 
32'd2000: dataIn1 = 32'd10; 
32'd2001: dataIn1 = 32'd39; 
32'd2002: dataIn1 = 32'd3; 
32'd2003: dataIn1 = 32'd14; 
32'd2004: dataIn1 = 32'd41; 
32'd2005: dataIn1 = 32'd16; 
32'd2006: dataIn1 = 32'd20; 
32'd2007: dataIn1 = 32'd26; 
32'd2008: dataIn1 = 32'd21; 
32'd2009: dataIn1 = 32'd14; 
32'd2010: dataIn1 = 32'd35; 
32'd2011: dataIn1 = 32'd45; 
32'd2012: dataIn1 = 32'd18; 
32'd2013: dataIn1 = 32'd42; 
32'd2014: dataIn1 = 32'd9; 
32'd2015: dataIn1 = 32'd60; 
32'd2016: dataIn1 = 32'd20; 
32'd2017: dataIn1 = 32'd62; 
32'd2018: dataIn1 = 32'd36; 
32'd2019: dataIn1 = 32'd63; 
32'd2020: dataIn1 = 32'd62; 
32'd2021: dataIn1 = 32'd61; 
32'd2022: dataIn1 = 32'd4; 
32'd2023: dataIn1 = 32'd26; 
32'd2024: dataIn1 = 32'd56; 
32'd2025: dataIn1 = 32'd41; 
32'd2026: dataIn1 = 32'd34; 
32'd2027: dataIn1 = 32'd15; 
32'd2028: dataIn1 = 32'd8; 
32'd2029: dataIn1 = 32'd14; 
32'd2030: dataIn1 = 32'd12; 
32'd2031: dataIn1 = 32'd3; 
32'd2032: dataIn1 = 32'd32; 
32'd2033: dataIn1 = 32'd13; 
32'd2034: dataIn1 = 32'd32; 
32'd2035: dataIn1 = 32'd42; 
32'd2036: dataIn1 = 32'd2; 
32'd2037: dataIn1 = 32'd50; 
32'd2038: dataIn1 = 32'd28; 
32'd2039: dataIn1 = 32'd50; 
32'd2040: dataIn1 = 32'd60; 
32'd2041: dataIn1 = 32'd57; 
32'd2042: dataIn1 = 32'd50; 
32'd2043: dataIn1 = 32'd36; 
32'd2044: dataIn1 = 32'd17; 
32'd2045: dataIn1 = 32'd41; 
32'd2046: dataIn1 = 32'd30; 
32'd2047: dataIn1 = 32'd47; 
32'd2048: dataIn1 = 32'd52; 
32'd2049: dataIn1 = 32'd14; 
32'd2050: dataIn1 = 32'd40; 
32'd2051: dataIn1 = 32'd63; 
32'd2052: dataIn1 = 32'd16; 
32'd2053: dataIn1 = 32'd9; 
32'd2054: dataIn1 = 32'd23; 
32'd2055: dataIn1 = 32'd16; 
32'd2056: dataIn1 = 32'd52; 
32'd2057: dataIn1 = 32'd41; 
32'd2058: dataIn1 = 32'd19; 
32'd2059: dataIn1 = 32'd31; 
32'd2060: dataIn1 = 32'd23; 
32'd2061: dataIn1 = 32'd8; 
32'd2062: dataIn1 = 32'd36; 
32'd2063: dataIn1 = 32'd2; 
32'd2064: dataIn1 = 32'd22; 
32'd2065: dataIn1 = 32'd38; 
32'd2066: dataIn1 = 32'd4; 
32'd2067: dataIn1 = 32'd15; 
32'd2068: dataIn1 = 32'd12; 
32'd2069: dataIn1 = 32'd4; 
32'd2070: dataIn1 = 32'd30; 
32'd2071: dataIn1 = 32'd30; 
32'd2072: dataIn1 = 32'd10; 
32'd2073: dataIn1 = 32'd2; 
32'd2074: dataIn1 = 32'd8; 
32'd2075: dataIn1 = 32'd13; 
32'd2076: dataIn1 = 32'd44; 
32'd2077: dataIn1 = 32'd34; 
32'd2078: dataIn1 = 32'd15; 
32'd2079: dataIn1 = 32'd56; 
32'd2080: dataIn1 = 32'd26; 
32'd2081: dataIn1 = 32'd56; 
32'd2082: dataIn1 = 32'd48; 
32'd2083: dataIn1 = 32'd59; 
32'd2084: dataIn1 = 32'd29; 
32'd2085: dataIn1 = 32'd48; 
32'd2086: dataIn1 = 32'd1; 
32'd2087: dataIn1 = 32'd38; 
32'd2088: dataIn1 = 32'd19; 
32'd2089: dataIn1 = 32'd32; 
32'd2090: dataIn1 = 32'd8; 
32'd2091: dataIn1 = 32'd13; 
32'd2092: dataIn1 = 32'd37; 
32'd2093: dataIn1 = 32'd25; 
32'd2094: dataIn1 = 32'd60; 
32'd2095: dataIn1 = 32'd30; 
32'd2096: dataIn1 = 32'd42; 
32'd2097: dataIn1 = 32'd22; 
32'd2098: dataIn1 = 32'd6; 
32'd2099: dataIn1 = 32'd25; 
32'd2100: dataIn1 = 32'd49; 
32'd2101: dataIn1 = 32'd3; 
32'd2102: dataIn1 = 32'd21; 
32'd2103: dataIn1 = 32'd7; 
32'd2104: dataIn1 = 32'd23; 
32'd2105: dataIn1 = 32'd7; 
32'd2106: dataIn1 = 32'd12; 
32'd2107: dataIn1 = 32'd50; 
32'd2108: dataIn1 = 32'd9; 
32'd2109: dataIn1 = 32'd22; 
32'd2110: dataIn1 = 32'd52; 
32'd2111: dataIn1 = 32'd63; 
32'd2112: dataIn1 = 32'd18; 
32'd2113: dataIn1 = 32'd40; 
32'd2114: dataIn1 = 32'd31; 
32'd2115: dataIn1 = 32'd53; 
32'd2116: dataIn1 = 32'd62; 
32'd2117: dataIn1 = 32'd22; 
32'd2118: dataIn1 = 32'd11; 
32'd2119: dataIn1 = 32'd62; 
32'd2120: dataIn1 = 32'd24; 
32'd2121: dataIn1 = 32'd26; 
32'd2122: dataIn1 = 32'd5; 
32'd2123: dataIn1 = 32'd47; 
32'd2124: dataIn1 = 32'd19; 
32'd2125: dataIn1 = 32'd27; 
32'd2126: dataIn1 = 32'd34; 
32'd2127: dataIn1 = 32'd11; 
32'd2128: dataIn1 = 32'd56; 
32'd2129: dataIn1 = 32'd31; 
32'd2130: dataIn1 = 32'd27; 
32'd2131: dataIn1 = 32'd57; 
32'd2132: dataIn1 = 32'd27; 
32'd2133: dataIn1 = 32'd59; 
32'd2134: dataIn1 = 32'd20; 
32'd2135: dataIn1 = 32'd34; 
32'd2136: dataIn1 = 32'd15; 
32'd2137: dataIn1 = 32'd12; 
32'd2138: dataIn1 = 32'd7; 
32'd2139: dataIn1 = 32'd8; 
32'd2140: dataIn1 = 32'd44; 
32'd2141: dataIn1 = 32'd20; 
32'd2142: dataIn1 = 32'd24; 
32'd2143: dataIn1 = 32'd41; 
32'd2144: dataIn1 = 32'd2; 
32'd2145: dataIn1 = 32'd30; 
32'd2146: dataIn1 = 32'd16; 
32'd2147: dataIn1 = 32'd33; 
32'd2148: dataIn1 = 32'd16; 
32'd2149: dataIn1 = 32'd27; 
32'd2150: dataIn1 = 32'd1; 
32'd2151: dataIn1 = 32'd36; 
32'd2152: dataIn1 = 32'd51; 
32'd2153: dataIn1 = 32'd2; 
32'd2154: dataIn1 = 32'd41; 
32'd2155: dataIn1 = 32'd36; 
32'd2156: dataIn1 = 32'd62; 
32'd2157: dataIn1 = 32'd57; 
32'd2158: dataIn1 = 32'd25; 
32'd2159: dataIn1 = 32'd57; 
32'd2160: dataIn1 = 32'd48; 
32'd2161: dataIn1 = 32'd17; 
32'd2162: dataIn1 = 32'd25; 
32'd2163: dataIn1 = 32'd39; 
32'd2164: dataIn1 = 32'd36; 
32'd2165: dataIn1 = 32'd16; 
32'd2166: dataIn1 = 32'd63; 
32'd2167: dataIn1 = 32'd16; 
32'd2168: dataIn1 = 32'd5; 
32'd2169: dataIn1 = 32'd58; 
32'd2170: dataIn1 = 32'd26; 
32'd2171: dataIn1 = 32'd1; 
32'd2172: dataIn1 = 32'd17; 
32'd2173: dataIn1 = 32'd39; 
32'd2174: dataIn1 = 32'd20; 
32'd2175: dataIn1 = 32'd58; 
32'd2176: dataIn1 = 32'd55; 
32'd2177: dataIn1 = 32'd17; 
32'd2178: dataIn1 = 32'd52; 
32'd2179: dataIn1 = 32'd44; 
32'd2180: dataIn1 = 32'd17; 
32'd2181: dataIn1 = 32'd61; 
32'd2182: dataIn1 = 32'd21; 
32'd2183: dataIn1 = 32'd20; 
32'd2184: dataIn1 = 32'd61; 
32'd2185: dataIn1 = 32'd56; 
32'd2186: dataIn1 = 32'd58; 
32'd2187: dataIn1 = 32'd57; 
32'd2188: dataIn1 = 32'd0; 
32'd2189: dataIn1 = 32'd35; 
32'd2190: dataIn1 = 32'd36; 
32'd2191: dataIn1 = 32'd31; 
32'd2192: dataIn1 = 32'd21; 
32'd2193: dataIn1 = 32'd2; 
32'd2194: dataIn1 = 32'd1; 
32'd2195: dataIn1 = 32'd27; 
32'd2196: dataIn1 = 32'd8; 
32'd2197: dataIn1 = 32'd58; 
32'd2198: dataIn1 = 32'd38; 
32'd2199: dataIn1 = 32'd43; 
32'd2200: dataIn1 = 32'd40; 
32'd2201: dataIn1 = 32'd58; 
32'd2202: dataIn1 = 32'd27; 
32'd2203: dataIn1 = 32'd37; 
32'd2204: dataIn1 = 32'd53; 
32'd2205: dataIn1 = 32'd38; 
32'd2206: dataIn1 = 32'd48; 
32'd2207: dataIn1 = 32'd13; 
32'd2208: dataIn1 = 32'd63; 
32'd2209: dataIn1 = 32'd21; 
32'd2210: dataIn1 = 32'd18; 
32'd2211: dataIn1 = 32'd6; 
32'd2212: dataIn1 = 32'd26; 
32'd2213: dataIn1 = 32'd63; 
32'd2214: dataIn1 = 32'd1; 
32'd2215: dataIn1 = 32'd0; 
32'd2216: dataIn1 = 32'd17; 
32'd2217: dataIn1 = 32'd63; 
32'd2218: dataIn1 = 32'd12; 
32'd2219: dataIn1 = 32'd20; 
32'd2220: dataIn1 = 32'd48; 
32'd2221: dataIn1 = 32'd10; 
32'd2222: dataIn1 = 32'd61; 
32'd2223: dataIn1 = 32'd24; 
32'd2224: dataIn1 = 32'd10; 
32'd2225: dataIn1 = 32'd4; 
32'd2226: dataIn1 = 32'd13; 
32'd2227: dataIn1 = 32'd15; 
32'd2228: dataIn1 = 32'd35; 
32'd2229: dataIn1 = 32'd57; 
32'd2230: dataIn1 = 32'd2; 
32'd2231: dataIn1 = 32'd34; 
32'd2232: dataIn1 = 32'd36; 
32'd2233: dataIn1 = 32'd56; 
32'd2234: dataIn1 = 32'd41; 
32'd2235: dataIn1 = 32'd3; 
32'd2236: dataIn1 = 32'd42; 
32'd2237: dataIn1 = 32'd63; 
32'd2238: dataIn1 = 32'd33; 
32'd2239: dataIn1 = 32'd63; 
32'd2240: dataIn1 = 32'd5; 
32'd2241: dataIn1 = 32'd23; 
32'd2242: dataIn1 = 32'd43; 
32'd2243: dataIn1 = 32'd24; 
32'd2244: dataIn1 = 32'd63; 
32'd2245: dataIn1 = 32'd51; 
32'd2246: dataIn1 = 32'd11; 
32'd2247: dataIn1 = 32'd6; 
32'd2248: dataIn1 = 32'd3; 
32'd2249: dataIn1 = 32'd4; 
32'd2250: dataIn1 = 32'd39; 
32'd2251: dataIn1 = 32'd6; 
32'd2252: dataIn1 = 32'd19; 
32'd2253: dataIn1 = 32'd9; 
32'd2254: dataIn1 = 32'd44; 
32'd2255: dataIn1 = 32'd6; 
32'd2256: dataIn1 = 32'd12; 
32'd2257: dataIn1 = 32'd13; 
32'd2258: dataIn1 = 32'd31; 
32'd2259: dataIn1 = 32'd52; 
32'd2260: dataIn1 = 32'd2; 
32'd2261: dataIn1 = 32'd57; 
32'd2262: dataIn1 = 32'd57; 
32'd2263: dataIn1 = 32'd2; 
32'd2264: dataIn1 = 32'd39; 
32'd2265: dataIn1 = 32'd31; 
32'd2266: dataIn1 = 32'd59; 
32'd2267: dataIn1 = 32'd62; 
32'd2268: dataIn1 = 32'd22; 
32'd2269: dataIn1 = 32'd62; 
32'd2270: dataIn1 = 32'd28; 
32'd2271: dataIn1 = 32'd48; 
32'd2272: dataIn1 = 32'd20; 
32'd2273: dataIn1 = 32'd60; 
32'd2274: dataIn1 = 32'd56; 
32'd2275: dataIn1 = 32'd17; 
32'd2276: dataIn1 = 32'd22; 
32'd2277: dataIn1 = 32'd11; 
32'd2278: dataIn1 = 32'd11; 
32'd2279: dataIn1 = 32'd19; 
32'd2280: dataIn1 = 32'd7; 
32'd2281: dataIn1 = 32'd24; 
32'd2282: dataIn1 = 32'd51; 
32'd2283: dataIn1 = 32'd50; 
32'd2284: dataIn1 = 32'd42; 
32'd2285: dataIn1 = 32'd19; 
32'd2286: dataIn1 = 32'd33; 
32'd2287: dataIn1 = 32'd9; 
32'd2288: dataIn1 = 32'd34; 
32'd2289: dataIn1 = 32'd52; 
32'd2290: dataIn1 = 32'd37; 
32'd2291: dataIn1 = 32'd61; 
32'd2292: dataIn1 = 32'd18; 
32'd2293: dataIn1 = 32'd20; 
32'd2294: dataIn1 = 32'd29; 
32'd2295: dataIn1 = 32'd49; 
32'd2296: dataIn1 = 32'd50; 
32'd2297: dataIn1 = 32'd31; 
32'd2298: dataIn1 = 32'd58; 
32'd2299: dataIn1 = 32'd2; 
32'd2300: dataIn1 = 32'd43; 
32'd2301: dataIn1 = 32'd33; 
32'd2302: dataIn1 = 32'd33; 
32'd2303: dataIn1 = 32'd4; 
32'd2304: dataIn1 = 32'd8; 
32'd2305: dataIn1 = 32'd15; 
32'd2306: dataIn1 = 32'd5; 
32'd2307: dataIn1 = 32'd55; 
32'd2308: dataIn1 = 32'd19; 
32'd2309: dataIn1 = 32'd21; 
32'd2310: dataIn1 = 32'd25; 
32'd2311: dataIn1 = 32'd29; 
32'd2312: dataIn1 = 32'd35; 
32'd2313: dataIn1 = 32'd27; 
32'd2314: dataIn1 = 32'd47; 
32'd2315: dataIn1 = 32'd27; 
32'd2316: dataIn1 = 32'd61; 
32'd2317: dataIn1 = 32'd56; 
32'd2318: dataIn1 = 32'd12; 
32'd2319: dataIn1 = 32'd48; 
32'd2320: dataIn1 = 32'd5; 
32'd2321: dataIn1 = 32'd22; 
32'd2322: dataIn1 = 32'd37; 
32'd2323: dataIn1 = 32'd11; 
32'd2324: dataIn1 = 32'd54; 
32'd2325: dataIn1 = 32'd39; 
32'd2326: dataIn1 = 32'd50; 
32'd2327: dataIn1 = 32'd22; 
32'd2328: dataIn1 = 32'd40; 
32'd2329: dataIn1 = 32'd32; 
32'd2330: dataIn1 = 32'd1; 
32'd2331: dataIn1 = 32'd34; 
32'd2332: dataIn1 = 32'd14; 
32'd2333: dataIn1 = 32'd11; 
32'd2334: dataIn1 = 32'd37; 
32'd2335: dataIn1 = 32'd62; 
32'd2336: dataIn1 = 32'd24; 
32'd2337: dataIn1 = 32'd36; 
32'd2338: dataIn1 = 32'd30; 
32'd2339: dataIn1 = 32'd10; 
32'd2340: dataIn1 = 32'd10; 
32'd2341: dataIn1 = 32'd41; 
32'd2342: dataIn1 = 32'd49; 
32'd2343: dataIn1 = 32'd32; 
32'd2344: dataIn1 = 32'd21; 
32'd2345: dataIn1 = 32'd61; 
32'd2346: dataIn1 = 32'd35; 
32'd2347: dataIn1 = 32'd38; 
32'd2348: dataIn1 = 32'd20; 
32'd2349: dataIn1 = 32'd49; 
32'd2350: dataIn1 = 32'd38; 
32'd2351: dataIn1 = 32'd16; 
32'd2352: dataIn1 = 32'd29; 
32'd2353: dataIn1 = 32'd45; 
32'd2354: dataIn1 = 32'd20; 
32'd2355: dataIn1 = 32'd34; 
32'd2356: dataIn1 = 32'd15; 
32'd2357: dataIn1 = 32'd62; 
32'd2358: dataIn1 = 32'd21; 
32'd2359: dataIn1 = 32'd15; 
32'd2360: dataIn1 = 32'd62; 
32'd2361: dataIn1 = 32'd5; 
32'd2362: dataIn1 = 32'd39; 
32'd2363: dataIn1 = 32'd29; 
32'd2364: dataIn1 = 32'd26; 
32'd2365: dataIn1 = 32'd28; 
32'd2366: dataIn1 = 32'd26; 
32'd2367: dataIn1 = 32'd50; 
32'd2368: dataIn1 = 32'd44; 
32'd2369: dataIn1 = 32'd48; 
32'd2370: dataIn1 = 32'd63; 
32'd2371: dataIn1 = 32'd23; 
32'd2372: dataIn1 = 32'd19; 
32'd2373: dataIn1 = 32'd63; 
32'd2374: dataIn1 = 32'd29; 
32'd2375: dataIn1 = 32'd17; 
32'd2376: dataIn1 = 32'd36; 
32'd2377: dataIn1 = 32'd50; 
32'd2378: dataIn1 = 32'd16; 
32'd2379: dataIn1 = 32'd55; 
32'd2380: dataIn1 = 32'd33; 
32'd2381: dataIn1 = 32'd40; 
32'd2382: dataIn1 = 32'd21; 
32'd2383: dataIn1 = 32'd56; 
32'd2384: dataIn1 = 32'd51; 
32'd2385: dataIn1 = 32'd44; 
32'd2386: dataIn1 = 32'd51; 
32'd2387: dataIn1 = 32'd40; 
32'd2388: dataIn1 = 32'd2; 
32'd2389: dataIn1 = 32'd11; 
32'd2390: dataIn1 = 32'd31; 
32'd2391: dataIn1 = 32'd29; 
32'd2392: dataIn1 = 32'd2; 
32'd2393: dataIn1 = 32'd42; 
32'd2394: dataIn1 = 32'd53; 
32'd2395: dataIn1 = 32'd26; 
32'd2396: dataIn1 = 32'd54; 
32'd2397: dataIn1 = 32'd25; 
32'd2398: dataIn1 = 32'd12; 
32'd2399: dataIn1 = 32'd44; 
32'd2400: dataIn1 = 32'd23; 
32'd2401: dataIn1 = 32'd21; 
32'd2402: dataIn1 = 32'd9; 
32'd2403: dataIn1 = 32'd52; 
32'd2404: dataIn1 = 32'd50; 
32'd2405: dataIn1 = 32'd37; 
32'd2406: dataIn1 = 32'd41; 
32'd2407: dataIn1 = 32'd60; 
32'd2408: dataIn1 = 32'd15; 
32'd2409: dataIn1 = 32'd42; 
32'd2410: dataIn1 = 32'd55; 
32'd2411: dataIn1 = 32'd31; 
32'd2412: dataIn1 = 32'd8; 
32'd2413: dataIn1 = 32'd18; 
32'd2414: dataIn1 = 32'd17; 
32'd2415: dataIn1 = 32'd29; 
32'd2416: dataIn1 = 32'd6; 
32'd2417: dataIn1 = 32'd48; 
32'd2418: dataIn1 = 32'd4; 
32'd2419: dataIn1 = 32'd59; 
32'd2420: dataIn1 = 32'd16; 
32'd2421: dataIn1 = 32'd16; 
32'd2422: dataIn1 = 32'd4; 
32'd2423: dataIn1 = 32'd2; 
32'd2424: dataIn1 = 32'd49; 
32'd2425: dataIn1 = 32'd28; 
32'd2426: dataIn1 = 32'd34; 
32'd2427: dataIn1 = 32'd34; 
32'd2428: dataIn1 = 32'd17; 
32'd2429: dataIn1 = 32'd34; 
32'd2430: dataIn1 = 32'd17; 
32'd2431: dataIn1 = 32'd45; 
32'd2432: dataIn1 = 32'd17; 
32'd2433: dataIn1 = 32'd5; 
32'd2434: dataIn1 = 32'd29; 
32'd2435: dataIn1 = 32'd19; 
32'd2436: dataIn1 = 32'd6; 
32'd2437: dataIn1 = 32'd14; 
32'd2438: dataIn1 = 32'd10; 
32'd2439: dataIn1 = 32'd56; 
32'd2440: dataIn1 = 32'd45; 
32'd2441: dataIn1 = 32'd11; 
32'd2442: dataIn1 = 32'd29; 
32'd2443: dataIn1 = 32'd11; 
32'd2444: dataIn1 = 32'd14; 
32'd2445: dataIn1 = 32'd62; 
32'd2446: dataIn1 = 32'd45; 
32'd2447: dataIn1 = 32'd22; 
32'd2448: dataIn1 = 32'd46; 
32'd2449: dataIn1 = 32'd43; 
32'd2450: dataIn1 = 32'd24; 
32'd2451: dataIn1 = 32'd17; 
32'd2452: dataIn1 = 32'd16; 
32'd2453: dataIn1 = 32'd61; 
32'd2454: dataIn1 = 32'd21; 
32'd2455: dataIn1 = 32'd51; 
32'd2456: dataIn1 = 32'd3; 
32'd2457: dataIn1 = 32'd29; 
32'd2458: dataIn1 = 32'd43; 
32'd2459: dataIn1 = 32'd18; 
32'd2460: dataIn1 = 32'd60; 
32'd2461: dataIn1 = 32'd43; 
32'd2462: dataIn1 = 32'd16; 
32'd2463: dataIn1 = 32'd12; 
32'd2464: dataIn1 = 32'd24; 
32'd2465: dataIn1 = 32'd62; 
32'd2466: dataIn1 = 32'd48; 
32'd2467: dataIn1 = 32'd63; 
32'd2468: dataIn1 = 32'd38; 
32'd2469: dataIn1 = 32'd14; 
32'd2470: dataIn1 = 32'd55; 
32'd2471: dataIn1 = 32'd5; 
32'd2472: dataIn1 = 32'd28; 
32'd2473: dataIn1 = 32'd35; 
32'd2474: dataIn1 = 32'd1; 
32'd2475: dataIn1 = 32'd19; 
32'd2476: dataIn1 = 32'd24; 
32'd2477: dataIn1 = 32'd28; 
32'd2478: dataIn1 = 32'd25; 
32'd2479: dataIn1 = 32'd44; 
32'd2480: dataIn1 = 32'd0; 
32'd2481: dataIn1 = 32'd55; 
32'd2482: dataIn1 = 32'd18; 
32'd2483: dataIn1 = 32'd22; 
32'd2484: dataIn1 = 32'd13; 
32'd2485: dataIn1 = 32'd2; 
32'd2486: dataIn1 = 32'd59; 
32'd2487: dataIn1 = 32'd2; 
32'd2488: dataIn1 = 32'd25; 
32'd2489: dataIn1 = 32'd10; 
32'd2490: dataIn1 = 32'd32; 
32'd2491: dataIn1 = 32'd55; 
32'd2492: dataIn1 = 32'd61; 
32'd2493: dataIn1 = 32'd3; 
32'd2494: dataIn1 = 32'd48; 
32'd2495: dataIn1 = 32'd44; 
32'd2496: dataIn1 = 32'd14; 
32'd2497: dataIn1 = 32'd3; 
32'd2498: dataIn1 = 32'd17; 
32'd2499: dataIn1 = 32'd60; 
32'd2500: dataIn1 = 32'd40; 
32'd2501: dataIn1 = 32'd24; 
32'd2502: dataIn1 = 32'd9; 
32'd2503: dataIn1 = 32'd40; 
32'd2504: dataIn1 = 32'd13; 
32'd2505: dataIn1 = 32'd35; 
32'd2506: dataIn1 = 32'd25; 
32'd2507: dataIn1 = 32'd47; 
32'd2508: dataIn1 = 32'd57; 
32'd2509: dataIn1 = 32'd31; 
32'd2510: dataIn1 = 32'd60; 
32'd2511: dataIn1 = 32'd21; 
32'd2512: dataIn1 = 32'd10; 
32'd2513: dataIn1 = 32'd36; 
32'd2514: dataIn1 = 32'd18; 
32'd2515: dataIn1 = 32'd21; 
32'd2516: dataIn1 = 32'd14; 
32'd2517: dataIn1 = 32'd59; 
32'd2518: dataIn1 = 32'd10; 
32'd2519: dataIn1 = 32'd45; 
32'd2520: dataIn1 = 32'd43; 
32'd2521: dataIn1 = 32'd4; 
32'd2522: dataIn1 = 32'd44; 
32'd2523: dataIn1 = 32'd9; 
32'd2524: dataIn1 = 32'd5; 
32'd2525: dataIn1 = 32'd50; 
32'd2526: dataIn1 = 32'd4; 
32'd2527: dataIn1 = 32'd28; 
32'd2528: dataIn1 = 32'd54; 
32'd2529: dataIn1 = 32'd7; 
32'd2530: dataIn1 = 32'd56; 
32'd2531: dataIn1 = 32'd28; 
32'd2532: dataIn1 = 32'd19; 
32'd2533: dataIn1 = 32'd21; 
32'd2534: dataIn1 = 32'd43; 
32'd2535: dataIn1 = 32'd25; 
32'd2536: dataIn1 = 32'd41; 
32'd2537: dataIn1 = 32'd18; 
32'd2538: dataIn1 = 32'd62; 
32'd2539: dataIn1 = 32'd18; 
32'd2540: dataIn1 = 32'd5; 
32'd2541: dataIn1 = 32'd10; 
32'd2542: dataIn1 = 32'd48; 
32'd2543: dataIn1 = 32'd45; 
32'd2544: dataIn1 = 32'd34; 
32'd2545: dataIn1 = 32'd32; 
32'd2546: dataIn1 = 32'd44; 
32'd2547: dataIn1 = 32'd61; 
32'd2548: dataIn1 = 32'd5; 
32'd2549: dataIn1 = 32'd51; 
32'd2550: dataIn1 = 32'd3; 
32'd2551: dataIn1 = 32'd32; 
32'd2552: dataIn1 = 32'd1; 
32'd2553: dataIn1 = 32'd44; 
32'd2554: dataIn1 = 32'd0; 
32'd2555: dataIn1 = 32'd14; 
32'd2556: dataIn1 = 32'd6; 
32'd2557: dataIn1 = 32'd62; 
32'd2558: dataIn1 = 32'd8; 
32'd2559: dataIn1 = 32'd55; 
32'd2560: dataIn1 = 32'd39; 
32'd2561: dataIn1 = 32'd5; 
32'd2562: dataIn1 = 32'd7; 
32'd2563: dataIn1 = 32'd57; 
32'd2564: dataIn1 = 32'd55; 
32'd2565: dataIn1 = 32'd24; 
32'd2566: dataIn1 = 32'd30; 
32'd2567: dataIn1 = 32'd35; 
32'd2568: dataIn1 = 32'd59; 
32'd2569: dataIn1 = 32'd9; 
32'd2570: dataIn1 = 32'd7; 
32'd2571: dataIn1 = 32'd29; 
32'd2572: dataIn1 = 32'd27; 
32'd2573: dataIn1 = 32'd11; 
32'd2574: dataIn1 = 32'd10; 
32'd2575: dataIn1 = 32'd54; 
32'd2576: dataIn1 = 32'd54; 
32'd2577: dataIn1 = 32'd28; 
32'd2578: dataIn1 = 32'd36; 
32'd2579: dataIn1 = 32'd30; 
32'd2580: dataIn1 = 32'd59; 
32'd2581: dataIn1 = 32'd51; 
32'd2582: dataIn1 = 32'd4; 
32'd2583: dataIn1 = 32'd45; 
32'd2584: dataIn1 = 32'd52; 
32'd2585: dataIn1 = 32'd30; 
32'd2586: dataIn1 = 32'd9; 
32'd2587: dataIn1 = 32'd37; 
32'd2588: dataIn1 = 32'd25; 
32'd2589: dataIn1 = 32'd49; 
32'd2590: dataIn1 = 32'd22; 
32'd2591: dataIn1 = 32'd39; 
32'd2592: dataIn1 = 32'd8; 
32'd2593: dataIn1 = 32'd30; 
32'd2594: dataIn1 = 32'd19; 
32'd2595: dataIn1 = 32'd17; 
32'd2596: dataIn1 = 32'd12; 
32'd2597: dataIn1 = 32'd32; 
32'd2598: dataIn1 = 32'd16; 
32'd2599: dataIn1 = 32'd34; 
32'd2600: dataIn1 = 32'd52; 
32'd2601: dataIn1 = 32'd17; 
32'd2602: dataIn1 = 32'd23; 
32'd2603: dataIn1 = 32'd49; 
32'd2604: dataIn1 = 32'd18; 
32'd2605: dataIn1 = 32'd20; 
32'd2606: dataIn1 = 32'd31; 
32'd2607: dataIn1 = 32'd15; 
32'd2608: dataIn1 = 32'd61; 
32'd2609: dataIn1 = 32'd48; 
32'd2610: dataIn1 = 32'd53; 
32'd2611: dataIn1 = 32'd47; 
32'd2612: dataIn1 = 32'd10; 
32'd2613: dataIn1 = 32'd3; 
32'd2614: dataIn1 = 32'd53; 
32'd2615: dataIn1 = 32'd21; 
32'd2616: dataIn1 = 32'd58; 
32'd2617: dataIn1 = 32'd11; 
32'd2618: dataIn1 = 32'd39; 
32'd2619: dataIn1 = 32'd61; 
32'd2620: dataIn1 = 32'd27; 
32'd2621: dataIn1 = 32'd17; 
32'd2622: dataIn1 = 32'd13; 
32'd2623: dataIn1 = 32'd14; 
32'd2624: dataIn1 = 32'd31; 
32'd2625: dataIn1 = 32'd30; 
32'd2626: dataIn1 = 32'd40; 
32'd2627: dataIn1 = 32'd63; 
32'd2628: dataIn1 = 32'd15; 
32'd2629: dataIn1 = 32'd23; 
32'd2630: dataIn1 = 32'd10; 
32'd2631: dataIn1 = 32'd25; 
32'd2632: dataIn1 = 32'd54; 
32'd2633: dataIn1 = 32'd56; 
32'd2634: dataIn1 = 32'd58; 
32'd2635: dataIn1 = 32'd26; 
32'd2636: dataIn1 = 32'd27; 
32'd2637: dataIn1 = 32'd12; 
32'd2638: dataIn1 = 32'd10; 
32'd2639: dataIn1 = 32'd15; 
32'd2640: dataIn1 = 32'd45; 
32'd2641: dataIn1 = 32'd56; 
32'd2642: dataIn1 = 32'd7; 
32'd2643: dataIn1 = 32'd59; 
32'd2644: dataIn1 = 32'd9; 
32'd2645: dataIn1 = 32'd46; 
32'd2646: dataIn1 = 32'd12; 
32'd2647: dataIn1 = 32'd34; 
32'd2648: dataIn1 = 32'd6; 
32'd2649: dataIn1 = 32'd48; 
32'd2650: dataIn1 = 32'd63; 
32'd2651: dataIn1 = 32'd8; 
32'd2652: dataIn1 = 32'd15; 
32'd2653: dataIn1 = 32'd3; 
32'd2654: dataIn1 = 32'd34; 
32'd2655: dataIn1 = 32'd60; 
32'd2656: dataIn1 = 32'd35; 
32'd2657: dataIn1 = 32'd1; 
32'd2658: dataIn1 = 32'd20; 
32'd2659: dataIn1 = 32'd55; 
32'd2660: dataIn1 = 32'd26; 
32'd2661: dataIn1 = 32'd47; 
32'd2662: dataIn1 = 32'd22; 
32'd2663: dataIn1 = 32'd5; 
32'd2664: dataIn1 = 32'd20; 
32'd2665: dataIn1 = 32'd8; 
32'd2666: dataIn1 = 32'd26; 
32'd2667: dataIn1 = 32'd18; 
32'd2668: dataIn1 = 32'd1; 
32'd2669: dataIn1 = 32'd45; 
32'd2670: dataIn1 = 32'd60; 
32'd2671: dataIn1 = 32'd41; 
32'd2672: dataIn1 = 32'd13; 
32'd2673: dataIn1 = 32'd42; 
32'd2674: dataIn1 = 32'd5; 
32'd2675: dataIn1 = 32'd5; 
32'd2676: dataIn1 = 32'd14; 
32'd2677: dataIn1 = 32'd13; 
32'd2678: dataIn1 = 32'd58; 
32'd2679: dataIn1 = 32'd6; 
32'd2680: dataIn1 = 32'd20; 
32'd2681: dataIn1 = 32'd16; 
32'd2682: dataIn1 = 32'd33; 
32'd2683: dataIn1 = 32'd6; 
32'd2684: dataIn1 = 32'd51; 
32'd2685: dataIn1 = 32'd11; 
32'd2686: dataIn1 = 32'd18; 
32'd2687: dataIn1 = 32'd14; 
32'd2688: dataIn1 = 32'd61; 
32'd2689: dataIn1 = 32'd55; 
32'd2690: dataIn1 = 32'd42; 
32'd2691: dataIn1 = 32'd1; 
32'd2692: dataIn1 = 32'd42; 
32'd2693: dataIn1 = 32'd11; 
32'd2694: dataIn1 = 32'd35; 
32'd2695: dataIn1 = 32'd29; 
32'd2696: dataIn1 = 32'd44; 
32'd2697: dataIn1 = 32'd44; 
32'd2698: dataIn1 = 32'd58; 
32'd2699: dataIn1 = 32'd21; 
32'd2700: dataIn1 = 32'd21; 
32'd2701: dataIn1 = 32'd62; 
32'd2702: dataIn1 = 32'd13; 
32'd2703: dataIn1 = 32'd52; 
32'd2704: dataIn1 = 32'd12; 
32'd2705: dataIn1 = 32'd15; 
32'd2706: dataIn1 = 32'd36; 
32'd2707: dataIn1 = 32'd53; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd60; 
32'd3: dataIn2 = 32'd86; 
32'd4: dataIn2 = 32'd24; 
32'd5: dataIn2 = 32'd33; 
32'd6: dataIn2 = 32'd9; 
32'd7: dataIn2 = 32'd19; 
32'd8: dataIn2 = 32'd4; 
32'd9: dataIn2 = 32'd42; 
32'd10: dataIn2 = 32'd16; 
32'd11: dataIn2 = 32'd90; 
32'd12: dataIn2 = 32'd56; 
32'd13: dataIn2 = 32'd26; 
32'd14: dataIn2 = 32'd62; 
32'd15: dataIn2 = 32'd49; 
32'd16: dataIn2 = 32'd97; 
32'd17: dataIn2 = 32'd0; 
32'd18: dataIn2 = 32'd47; 
32'd19: dataIn2 = 32'd4; 
32'd20: dataIn2 = 32'd76; 
32'd21: dataIn2 = 32'd67; 
32'd22: dataIn2 = 32'd100; 
32'd23: dataIn2 = 32'd30; 
32'd24: dataIn2 = 32'd86; 
32'd25: dataIn2 = 32'd42; 
32'd26: dataIn2 = 32'd4; 
32'd27: dataIn2 = 32'd95; 
32'd28: dataIn2 = 32'd36; 
32'd29: dataIn2 = 32'd56; 
32'd30: dataIn2 = 32'd25; 
32'd31: dataIn2 = 32'd52; 
32'd32: dataIn2 = 32'd47; 
32'd33: dataIn2 = 32'd62; 
32'd34: dataIn2 = 32'd49; 
32'd35: dataIn2 = 32'd9; 
32'd36: dataIn2 = 32'd62; 
32'd37: dataIn2 = 32'd95; 
32'd38: dataIn2 = 32'd3; 
32'd39: dataIn2 = 32'd29; 
32'd40: dataIn2 = 32'd27; 
32'd41: dataIn2 = 32'd54; 
32'd42: dataIn2 = 32'd52; 
32'd43: dataIn2 = 32'd96; 
32'd44: dataIn2 = 32'd24; 
32'd45: dataIn2 = 32'd73; 
32'd46: dataIn2 = 32'd56; 
32'd47: dataIn2 = 32'd30; 
32'd48: dataIn2 = 32'd13; 
32'd49: dataIn2 = 32'd38; 
32'd50: dataIn2 = 32'd60; 
32'd51: dataIn2 = 32'd47; 
32'd52: dataIn2 = 32'd3; 
32'd53: dataIn2 = 32'd4; 
32'd54: dataIn2 = 32'd85; 
32'd55: dataIn2 = 32'd53; 
32'd56: dataIn2 = 32'd40; 
32'd57: dataIn2 = 32'd93; 
32'd58: dataIn2 = 32'd44; 
32'd59: dataIn2 = 32'd83; 
32'd60: dataIn2 = 32'd100; 
32'd61: dataIn2 = 32'd34; 
32'd62: dataIn2 = 32'd6; 
32'd63: dataIn2 = 32'd80; 
32'd64: dataIn2 = 32'd45; 
32'd65: dataIn2 = 32'd42; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht1_64_50.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
