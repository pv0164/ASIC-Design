//64x64 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 1638 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd330 ; 
  wdata_col_base = 32'd19680 ; 
  row_base = 32'd213180 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #179000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd213180: dataIn1 = 32'd0
; 
32'd213181: dataIn1 = 32'd25
; 
32'd213182: dataIn1 = 32'd50
; 
32'd213183: dataIn1 = 32'd81
; 
32'd213184: dataIn1 = 32'd106
; 
32'd213185: dataIn1 = 32'd130
; 
32'd213186: dataIn1 = 32'd149
; 
32'd213187: dataIn1 = 32'd182
; 
32'd213188: dataIn1 = 32'd206
; 
32'd213189: dataIn1 = 32'd233
; 
32'd213190: dataIn1 = 32'd258
; 
32'd213191: dataIn1 = 32'd279
; 
32'd213192: dataIn1 = 32'd306
; 
32'd213193: dataIn1 = 32'd337
; 
32'd213194: dataIn1 = 32'd362
; 
32'd213195: dataIn1 = 32'd394
; 
32'd213196: dataIn1 = 32'd417
; 
32'd213197: dataIn1 = 32'd437
; 
32'd213198: dataIn1 = 32'd463
; 
32'd213199: dataIn1 = 32'd487
; 
32'd213200: dataIn1 = 32'd511
; 
32'd213201: dataIn1 = 32'd537
; 
32'd213202: dataIn1 = 32'd564
; 
32'd213203: dataIn1 = 32'd590
; 
32'd213204: dataIn1 = 32'd613
; 
32'd213205: dataIn1 = 32'd639
; 
32'd213206: dataIn1 = 32'd664
; 
32'd213207: dataIn1 = 32'd682
; 
32'd213208: dataIn1 = 32'd706
; 
32'd213209: dataIn1 = 32'd726
; 
32'd213210: dataIn1 = 32'd750
; 
32'd213211: dataIn1 = 32'd774
; 
32'd213212: dataIn1 = 32'd797
; 
32'd213213: dataIn1 = 32'd827
; 
32'd213214: dataIn1 = 32'd856
; 
32'd213215: dataIn1 = 32'd878
; 
32'd213216: dataIn1 = 32'd901
; 
32'd213217: dataIn1 = 32'd920
; 
32'd213218: dataIn1 = 32'd947
; 
32'd213219: dataIn1 = 32'd972
; 
32'd213220: dataIn1 = 32'd995
; 
32'd213221: dataIn1 = 32'd1014
; 
32'd213222: dataIn1 = 32'd1032
; 
32'd213223: dataIn1 = 32'd1056
; 
32'd213224: dataIn1 = 32'd1080
; 
32'd213225: dataIn1 = 32'd1106
; 
32'd213226: dataIn1 = 32'd1131
; 
32'd213227: dataIn1 = 32'd1152
; 
32'd213228: dataIn1 = 32'd1176
; 
32'd213229: dataIn1 = 32'd1194
; 
32'd213230: dataIn1 = 32'd1215
; 
32'd213231: dataIn1 = 32'd1236
; 
32'd213232: dataIn1 = 32'd1265
; 
32'd213233: dataIn1 = 32'd1293
; 
32'd213234: dataIn1 = 32'd1322
; 
32'd213235: dataIn1 = 32'd1346
; 
32'd213236: dataIn1 = 32'd1377
; 
32'd213237: dataIn1 = 32'd1405
; 
32'd213238: dataIn1 = 32'd1431
; 
32'd213239: dataIn1 = 32'd1457
; 
32'd213240: dataIn1 = 32'd1481
; 
32'd213241: dataIn1 = 32'd1503
; 
32'd213242: dataIn1 = 32'd1522
; 
32'd213243: dataIn1 = 32'd1543
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd19680: dataIn1 = 32'd0
; 
32'd19681: dataIn1 = 32'd25
; 
32'd19682: dataIn1 = 32'd50
; 
32'd19683: dataIn1 = 32'd81
; 
32'd19684: dataIn1 = 32'd106
; 
32'd19685: dataIn1 = 32'd130
; 
32'd19686: dataIn1 = 32'd149
; 
32'd19687: dataIn1 = 32'd182
; 
32'd19688: dataIn1 = 32'd206
; 
32'd19689: dataIn1 = 32'd233
; 
32'd19690: dataIn1 = 32'd258
; 
32'd19691: dataIn1 = 32'd279
; 
32'd19692: dataIn1 = 32'd306
; 
32'd19693: dataIn1 = 32'd337
; 
32'd19694: dataIn1 = 32'd362
; 
32'd19695: dataIn1 = 32'd394
; 
32'd19696: dataIn1 = 32'd417
; 
32'd19697: dataIn1 = 32'd437
; 
32'd19698: dataIn1 = 32'd463
; 
32'd19699: dataIn1 = 32'd487
; 
32'd19700: dataIn1 = 32'd511
; 
32'd19701: dataIn1 = 32'd537
; 
32'd19702: dataIn1 = 32'd564
; 
32'd19703: dataIn1 = 32'd590
; 
32'd19704: dataIn1 = 32'd613
; 
32'd19705: dataIn1 = 32'd639
; 
32'd19706: dataIn1 = 32'd664
; 
32'd19707: dataIn1 = 32'd682
; 
32'd19708: dataIn1 = 32'd706
; 
32'd19709: dataIn1 = 32'd726
; 
32'd19710: dataIn1 = 32'd750
; 
32'd19711: dataIn1 = 32'd774
; 
32'd19712: dataIn1 = 32'd797
; 
32'd19713: dataIn1 = 32'd827
; 
32'd19714: dataIn1 = 32'd856
; 
32'd19715: dataIn1 = 32'd878
; 
32'd19716: dataIn1 = 32'd901
; 
32'd19717: dataIn1 = 32'd920
; 
32'd19718: dataIn1 = 32'd947
; 
32'd19719: dataIn1 = 32'd972
; 
32'd19720: dataIn1 = 32'd995
; 
32'd19721: dataIn1 = 32'd1014
; 
32'd19722: dataIn1 = 32'd1032
; 
32'd19723: dataIn1 = 32'd1056
; 
32'd19724: dataIn1 = 32'd1080
; 
32'd19725: dataIn1 = 32'd1106
; 
32'd19726: dataIn1 = 32'd1131
; 
32'd19727: dataIn1 = 32'd1152
; 
32'd19728: dataIn1 = 32'd1176
; 
32'd19729: dataIn1 = 32'd1194
; 
32'd19730: dataIn1 = 32'd1215
; 
32'd19731: dataIn1 = 32'd1236
; 
32'd19732: dataIn1 = 32'd1265
; 
32'd19733: dataIn1 = 32'd1293
; 
32'd19734: dataIn1 = 32'd1322
; 
32'd19735: dataIn1 = 32'd1346
; 
32'd19736: dataIn1 = 32'd1377
; 
32'd19737: dataIn1 = 32'd1405
; 
32'd19738: dataIn1 = 32'd1431
; 
32'd19739: dataIn1 = 32'd1457
; 
32'd19740: dataIn1 = 32'd1481
; 
32'd19741: dataIn1 = 32'd1503
; 
32'd19742: dataIn1 = 32'd1522
; 
32'd19743: dataIn1 = 32'd1543
; 
32'd19744: dataIn1 = 32'd1557
; 
32'd19745: dataIn1 = 32'd2
; 
32'd19746: dataIn1 = 32'd3
; 
32'd19747: dataIn1 = 32'd5
; 
32'd19748: dataIn1 = 32'd10
; 
32'd19749: dataIn1 = 32'd12
; 
32'd19750: dataIn1 = 32'd17
; 
32'd19751: dataIn1 = 32'd18
; 
32'd19752: dataIn1 = 32'd20
; 
32'd19753: dataIn1 = 32'd27
; 
32'd19754: dataIn1 = 32'd29
; 
32'd19755: dataIn1 = 32'd30
; 
32'd19756: dataIn1 = 32'd31
; 
32'd19757: dataIn1 = 32'd32
; 
32'd19758: dataIn1 = 32'd33
; 
32'd19759: dataIn1 = 32'd35
; 
32'd19760: dataIn1 = 32'd37
; 
32'd19761: dataIn1 = 32'd41
; 
32'd19762: dataIn1 = 32'd42
; 
32'd19763: dataIn1 = 32'd46
; 
32'd19764: dataIn1 = 32'd47
; 
32'd19765: dataIn1 = 32'd49
; 
32'd19766: dataIn1 = 32'd54
; 
32'd19767: dataIn1 = 32'd58
; 
32'd19768: dataIn1 = 32'd59
; 
32'd19769: dataIn1 = 32'd61
; 
32'd19770: dataIn1 = 32'd6
; 
32'd19771: dataIn1 = 32'd7
; 
32'd19772: dataIn1 = 32'd8
; 
32'd19773: dataIn1 = 32'd9
; 
32'd19774: dataIn1 = 32'd13
; 
32'd19775: dataIn1 = 32'd15
; 
32'd19776: dataIn1 = 32'd20
; 
32'd19777: dataIn1 = 32'd21
; 
32'd19778: dataIn1 = 32'd22
; 
32'd19779: dataIn1 = 32'd23
; 
32'd19780: dataIn1 = 32'd24
; 
32'd19781: dataIn1 = 32'd29
; 
32'd19782: dataIn1 = 32'd31
; 
32'd19783: dataIn1 = 32'd32
; 
32'd19784: dataIn1 = 32'd34
; 
32'd19785: dataIn1 = 32'd36
; 
32'd19786: dataIn1 = 32'd38
; 
32'd19787: dataIn1 = 32'd39
; 
32'd19788: dataIn1 = 32'd41
; 
32'd19789: dataIn1 = 32'd42
; 
32'd19790: dataIn1 = 32'd50
; 
32'd19791: dataIn1 = 32'd52
; 
32'd19792: dataIn1 = 32'd57
; 
32'd19793: dataIn1 = 32'd60
; 
32'd19794: dataIn1 = 32'd63
; 
32'd19795: dataIn1 = 32'd0
; 
32'd19796: dataIn1 = 32'd1
; 
32'd19797: dataIn1 = 32'd2
; 
32'd19798: dataIn1 = 32'd3
; 
32'd19799: dataIn1 = 32'd4
; 
32'd19800: dataIn1 = 32'd8
; 
32'd19801: dataIn1 = 32'd9
; 
32'd19802: dataIn1 = 32'd12
; 
32'd19803: dataIn1 = 32'd13
; 
32'd19804: dataIn1 = 32'd14
; 
32'd19805: dataIn1 = 32'd18
; 
32'd19806: dataIn1 = 32'd19
; 
32'd19807: dataIn1 = 32'd21
; 
32'd19808: dataIn1 = 32'd24
; 
32'd19809: dataIn1 = 32'd25
; 
32'd19810: dataIn1 = 32'd26
; 
32'd19811: dataIn1 = 32'd28
; 
32'd19812: dataIn1 = 32'd29
; 
32'd19813: dataIn1 = 32'd30
; 
32'd19814: dataIn1 = 32'd34
; 
32'd19815: dataIn1 = 32'd36
; 
32'd19816: dataIn1 = 32'd38
; 
32'd19817: dataIn1 = 32'd40
; 
32'd19818: dataIn1 = 32'd46
; 
32'd19819: dataIn1 = 32'd52
; 
32'd19820: dataIn1 = 32'd53
; 
32'd19821: dataIn1 = 32'd54
; 
32'd19822: dataIn1 = 32'd56
; 
32'd19823: dataIn1 = 32'd58
; 
32'd19824: dataIn1 = 32'd60
; 
32'd19825: dataIn1 = 32'd61
; 
32'd19826: dataIn1 = 32'd1
; 
32'd19827: dataIn1 = 32'd4
; 
32'd19828: dataIn1 = 32'd6
; 
32'd19829: dataIn1 = 32'd7
; 
32'd19830: dataIn1 = 32'd8
; 
32'd19831: dataIn1 = 32'd10
; 
32'd19832: dataIn1 = 32'd11
; 
32'd19833: dataIn1 = 32'd13
; 
32'd19834: dataIn1 = 32'd18
; 
32'd19835: dataIn1 = 32'd24
; 
32'd19836: dataIn1 = 32'd29
; 
32'd19837: dataIn1 = 32'd30
; 
32'd19838: dataIn1 = 32'd31
; 
32'd19839: dataIn1 = 32'd33
; 
32'd19840: dataIn1 = 32'd39
; 
32'd19841: dataIn1 = 32'd40
; 
32'd19842: dataIn1 = 32'd42
; 
32'd19843: dataIn1 = 32'd43
; 
32'd19844: dataIn1 = 32'd45
; 
32'd19845: dataIn1 = 32'd47
; 
32'd19846: dataIn1 = 32'd51
; 
32'd19847: dataIn1 = 32'd53
; 
32'd19848: dataIn1 = 32'd58
; 
32'd19849: dataIn1 = 32'd60
; 
32'd19850: dataIn1 = 32'd63
; 
32'd19851: dataIn1 = 32'd0
; 
32'd19852: dataIn1 = 32'd3
; 
32'd19853: dataIn1 = 32'd5
; 
32'd19854: dataIn1 = 32'd17
; 
32'd19855: dataIn1 = 32'd18
; 
32'd19856: dataIn1 = 32'd19
; 
32'd19857: dataIn1 = 32'd21
; 
32'd19858: dataIn1 = 32'd24
; 
32'd19859: dataIn1 = 32'd26
; 
32'd19860: dataIn1 = 32'd28
; 
32'd19861: dataIn1 = 32'd31
; 
32'd19862: dataIn1 = 32'd39
; 
32'd19863: dataIn1 = 32'd40
; 
32'd19864: dataIn1 = 32'd43
; 
32'd19865: dataIn1 = 32'd44
; 
32'd19866: dataIn1 = 32'd45
; 
32'd19867: dataIn1 = 32'd50
; 
32'd19868: dataIn1 = 32'd52
; 
32'd19869: dataIn1 = 32'd54
; 
32'd19870: dataIn1 = 32'd56
; 
32'd19871: dataIn1 = 32'd59
; 
32'd19872: dataIn1 = 32'd60
; 
32'd19873: dataIn1 = 32'd61
; 
32'd19874: dataIn1 = 32'd63
; 
32'd19875: dataIn1 = 32'd0
; 
32'd19876: dataIn1 = 32'd2
; 
32'd19877: dataIn1 = 32'd10
; 
32'd19878: dataIn1 = 32'd11
; 
32'd19879: dataIn1 = 32'd16
; 
32'd19880: dataIn1 = 32'd18
; 
32'd19881: dataIn1 = 32'd19
; 
32'd19882: dataIn1 = 32'd21
; 
32'd19883: dataIn1 = 32'd22
; 
32'd19884: dataIn1 = 32'd23
; 
32'd19885: dataIn1 = 32'd35
; 
32'd19886: dataIn1 = 32'd40
; 
32'd19887: dataIn1 = 32'd41
; 
32'd19888: dataIn1 = 32'd46
; 
32'd19889: dataIn1 = 32'd48
; 
32'd19890: dataIn1 = 32'd49
; 
32'd19891: dataIn1 = 32'd50
; 
32'd19892: dataIn1 = 32'd54
; 
32'd19893: dataIn1 = 32'd58
; 
32'd19894: dataIn1 = 32'd2
; 
32'd19895: dataIn1 = 32'd3
; 
32'd19896: dataIn1 = 32'd4
; 
32'd19897: dataIn1 = 32'd6
; 
32'd19898: dataIn1 = 32'd7
; 
32'd19899: dataIn1 = 32'd10
; 
32'd19900: dataIn1 = 32'd11
; 
32'd19901: dataIn1 = 32'd13
; 
32'd19902: dataIn1 = 32'd15
; 
32'd19903: dataIn1 = 32'd16
; 
32'd19904: dataIn1 = 32'd17
; 
32'd19905: dataIn1 = 32'd18
; 
32'd19906: dataIn1 = 32'd20
; 
32'd19907: dataIn1 = 32'd21
; 
32'd19908: dataIn1 = 32'd22
; 
32'd19909: dataIn1 = 32'd24
; 
32'd19910: dataIn1 = 32'd25
; 
32'd19911: dataIn1 = 32'd27
; 
32'd19912: dataIn1 = 32'd29
; 
32'd19913: dataIn1 = 32'd30
; 
32'd19914: dataIn1 = 32'd31
; 
32'd19915: dataIn1 = 32'd34
; 
32'd19916: dataIn1 = 32'd35
; 
32'd19917: dataIn1 = 32'd40
; 
32'd19918: dataIn1 = 32'd43
; 
32'd19919: dataIn1 = 32'd46
; 
32'd19920: dataIn1 = 32'd47
; 
32'd19921: dataIn1 = 32'd48
; 
32'd19922: dataIn1 = 32'd49
; 
32'd19923: dataIn1 = 32'd55
; 
32'd19924: dataIn1 = 32'd56
; 
32'd19925: dataIn1 = 32'd57
; 
32'd19926: dataIn1 = 32'd62
; 
32'd19927: dataIn1 = 32'd1
; 
32'd19928: dataIn1 = 32'd5
; 
32'd19929: dataIn1 = 32'd7
; 
32'd19930: dataIn1 = 32'd10
; 
32'd19931: dataIn1 = 32'd14
; 
32'd19932: dataIn1 = 32'd15
; 
32'd19933: dataIn1 = 32'd23
; 
32'd19934: dataIn1 = 32'd25
; 
32'd19935: dataIn1 = 32'd27
; 
32'd19936: dataIn1 = 32'd28
; 
32'd19937: dataIn1 = 32'd30
; 
32'd19938: dataIn1 = 32'd31
; 
32'd19939: dataIn1 = 32'd32
; 
32'd19940: dataIn1 = 32'd34
; 
32'd19941: dataIn1 = 32'd36
; 
32'd19942: dataIn1 = 32'd37
; 
32'd19943: dataIn1 = 32'd39
; 
32'd19944: dataIn1 = 32'd41
; 
32'd19945: dataIn1 = 32'd42
; 
32'd19946: dataIn1 = 32'd44
; 
32'd19947: dataIn1 = 32'd48
; 
32'd19948: dataIn1 = 32'd50
; 
32'd19949: dataIn1 = 32'd56
; 
32'd19950: dataIn1 = 32'd62
; 
32'd19951: dataIn1 = 32'd2
; 
32'd19952: dataIn1 = 32'd6
; 
32'd19953: dataIn1 = 32'd9
; 
32'd19954: dataIn1 = 32'd13
; 
32'd19955: dataIn1 = 32'd25
; 
32'd19956: dataIn1 = 32'd26
; 
32'd19957: dataIn1 = 32'd32
; 
32'd19958: dataIn1 = 32'd33
; 
32'd19959: dataIn1 = 32'd34
; 
32'd19960: dataIn1 = 32'd36
; 
32'd19961: dataIn1 = 32'd37
; 
32'd19962: dataIn1 = 32'd39
; 
32'd19963: dataIn1 = 32'd40
; 
32'd19964: dataIn1 = 32'd41
; 
32'd19965: dataIn1 = 32'd42
; 
32'd19966: dataIn1 = 32'd43
; 
32'd19967: dataIn1 = 32'd45
; 
32'd19968: dataIn1 = 32'd46
; 
32'd19969: dataIn1 = 32'd47
; 
32'd19970: dataIn1 = 32'd48
; 
32'd19971: dataIn1 = 32'd54
; 
32'd19972: dataIn1 = 32'd55
; 
32'd19973: dataIn1 = 32'd56
; 
32'd19974: dataIn1 = 32'd57
; 
32'd19975: dataIn1 = 32'd58
; 
32'd19976: dataIn1 = 32'd60
; 
32'd19977: dataIn1 = 32'd63
; 
32'd19978: dataIn1 = 32'd3
; 
32'd19979: dataIn1 = 32'd5
; 
32'd19980: dataIn1 = 32'd6
; 
32'd19981: dataIn1 = 32'd8
; 
32'd19982: dataIn1 = 32'd10
; 
32'd19983: dataIn1 = 32'd12
; 
32'd19984: dataIn1 = 32'd15
; 
32'd19985: dataIn1 = 32'd16
; 
32'd19986: dataIn1 = 32'd19
; 
32'd19987: dataIn1 = 32'd25
; 
32'd19988: dataIn1 = 32'd34
; 
32'd19989: dataIn1 = 32'd36
; 
32'd19990: dataIn1 = 32'd37
; 
32'd19991: dataIn1 = 32'd38
; 
32'd19992: dataIn1 = 32'd39
; 
32'd19993: dataIn1 = 32'd40
; 
32'd19994: dataIn1 = 32'd43
; 
32'd19995: dataIn1 = 32'd47
; 
32'd19996: dataIn1 = 32'd48
; 
32'd19997: dataIn1 = 32'd49
; 
32'd19998: dataIn1 = 32'd50
; 
32'd19999: dataIn1 = 32'd51
; 
32'd20000: dataIn1 = 32'd53
; 
32'd20001: dataIn1 = 32'd55
; 
32'd20002: dataIn1 = 32'd57
; 
32'd20003: dataIn1 = 32'd0
; 
32'd20004: dataIn1 = 32'd1
; 
32'd20005: dataIn1 = 32'd2
; 
32'd20006: dataIn1 = 32'd7
; 
32'd20007: dataIn1 = 32'd16
; 
32'd20008: dataIn1 = 32'd17
; 
32'd20009: dataIn1 = 32'd18
; 
32'd20010: dataIn1 = 32'd22
; 
32'd20011: dataIn1 = 32'd23
; 
32'd20012: dataIn1 = 32'd24
; 
32'd20013: dataIn1 = 32'd27
; 
32'd20014: dataIn1 = 32'd34
; 
32'd20015: dataIn1 = 32'd36
; 
32'd20016: dataIn1 = 32'd37
; 
32'd20017: dataIn1 = 32'd38
; 
32'd20018: dataIn1 = 32'd46
; 
32'd20019: dataIn1 = 32'd50
; 
32'd20020: dataIn1 = 32'd51
; 
32'd20021: dataIn1 = 32'd55
; 
32'd20022: dataIn1 = 32'd56
; 
32'd20023: dataIn1 = 32'd60
; 
32'd20024: dataIn1 = 32'd1
; 
32'd20025: dataIn1 = 32'd2
; 
32'd20026: dataIn1 = 32'd3
; 
32'd20027: dataIn1 = 32'd5
; 
32'd20028: dataIn1 = 32'd7
; 
32'd20029: dataIn1 = 32'd8
; 
32'd20030: dataIn1 = 32'd10
; 
32'd20031: dataIn1 = 32'd11
; 
32'd20032: dataIn1 = 32'd14
; 
32'd20033: dataIn1 = 32'd15
; 
32'd20034: dataIn1 = 32'd16
; 
32'd20035: dataIn1 = 32'd18
; 
32'd20036: dataIn1 = 32'd19
; 
32'd20037: dataIn1 = 32'd20
; 
32'd20038: dataIn1 = 32'd21
; 
32'd20039: dataIn1 = 32'd22
; 
32'd20040: dataIn1 = 32'd26
; 
32'd20041: dataIn1 = 32'd30
; 
32'd20042: dataIn1 = 32'd33
; 
32'd20043: dataIn1 = 32'd40
; 
32'd20044: dataIn1 = 32'd46
; 
32'd20045: dataIn1 = 32'd47
; 
32'd20046: dataIn1 = 32'd48
; 
32'd20047: dataIn1 = 32'd50
; 
32'd20048: dataIn1 = 32'd53
; 
32'd20049: dataIn1 = 32'd56
; 
32'd20050: dataIn1 = 32'd58
; 
32'd20051: dataIn1 = 32'd0
; 
32'd20052: dataIn1 = 32'd2
; 
32'd20053: dataIn1 = 32'd6
; 
32'd20054: dataIn1 = 32'd8
; 
32'd20055: dataIn1 = 32'd12
; 
32'd20056: dataIn1 = 32'd13
; 
32'd20057: dataIn1 = 32'd20
; 
32'd20058: dataIn1 = 32'd21
; 
32'd20059: dataIn1 = 32'd23
; 
32'd20060: dataIn1 = 32'd27
; 
32'd20061: dataIn1 = 32'd28
; 
32'd20062: dataIn1 = 32'd29
; 
32'd20063: dataIn1 = 32'd30
; 
32'd20064: dataIn1 = 32'd31
; 
32'd20065: dataIn1 = 32'd33
; 
32'd20066: dataIn1 = 32'd34
; 
32'd20067: dataIn1 = 32'd36
; 
32'd20068: dataIn1 = 32'd38
; 
32'd20069: dataIn1 = 32'd39
; 
32'd20070: dataIn1 = 32'd41
; 
32'd20071: dataIn1 = 32'd42
; 
32'd20072: dataIn1 = 32'd45
; 
32'd20073: dataIn1 = 32'd46
; 
32'd20074: dataIn1 = 32'd47
; 
32'd20075: dataIn1 = 32'd49
; 
32'd20076: dataIn1 = 32'd51
; 
32'd20077: dataIn1 = 32'd53
; 
32'd20078: dataIn1 = 32'd57
; 
32'd20079: dataIn1 = 32'd59
; 
32'd20080: dataIn1 = 32'd60
; 
32'd20081: dataIn1 = 32'd61
; 
32'd20082: dataIn1 = 32'd2
; 
32'd20083: dataIn1 = 32'd11
; 
32'd20084: dataIn1 = 32'd12
; 
32'd20085: dataIn1 = 32'd14
; 
32'd20086: dataIn1 = 32'd15
; 
32'd20087: dataIn1 = 32'd16
; 
32'd20088: dataIn1 = 32'd17
; 
32'd20089: dataIn1 = 32'd18
; 
32'd20090: dataIn1 = 32'd20
; 
32'd20091: dataIn1 = 32'd21
; 
32'd20092: dataIn1 = 32'd25
; 
32'd20093: dataIn1 = 32'd27
; 
32'd20094: dataIn1 = 32'd28
; 
32'd20095: dataIn1 = 32'd33
; 
32'd20096: dataIn1 = 32'd34
; 
32'd20097: dataIn1 = 32'd36
; 
32'd20098: dataIn1 = 32'd43
; 
32'd20099: dataIn1 = 32'd44
; 
32'd20100: dataIn1 = 32'd49
; 
32'd20101: dataIn1 = 32'd50
; 
32'd20102: dataIn1 = 32'd51
; 
32'd20103: dataIn1 = 32'd59
; 
32'd20104: dataIn1 = 32'd60
; 
32'd20105: dataIn1 = 32'd61
; 
32'd20106: dataIn1 = 32'd62
; 
32'd20107: dataIn1 = 32'd1
; 
32'd20108: dataIn1 = 32'd3
; 
32'd20109: dataIn1 = 32'd10
; 
32'd20110: dataIn1 = 32'd17
; 
32'd20111: dataIn1 = 32'd18
; 
32'd20112: dataIn1 = 32'd21
; 
32'd20113: dataIn1 = 32'd22
; 
32'd20114: dataIn1 = 32'd23
; 
32'd20115: dataIn1 = 32'd26
; 
32'd20116: dataIn1 = 32'd30
; 
32'd20117: dataIn1 = 32'd32
; 
32'd20118: dataIn1 = 32'd33
; 
32'd20119: dataIn1 = 32'd34
; 
32'd20120: dataIn1 = 32'd35
; 
32'd20121: dataIn1 = 32'd38
; 
32'd20122: dataIn1 = 32'd39
; 
32'd20123: dataIn1 = 32'd42
; 
32'd20124: dataIn1 = 32'd43
; 
32'd20125: dataIn1 = 32'd44
; 
32'd20126: dataIn1 = 32'd45
; 
32'd20127: dataIn1 = 32'd46
; 
32'd20128: dataIn1 = 32'd47
; 
32'd20129: dataIn1 = 32'd48
; 
32'd20130: dataIn1 = 32'd51
; 
32'd20131: dataIn1 = 32'd54
; 
32'd20132: dataIn1 = 32'd55
; 
32'd20133: dataIn1 = 32'd56
; 
32'd20134: dataIn1 = 32'd58
; 
32'd20135: dataIn1 = 32'd59
; 
32'd20136: dataIn1 = 32'd60
; 
32'd20137: dataIn1 = 32'd62
; 
32'd20138: dataIn1 = 32'd63
; 
32'd20139: dataIn1 = 32'd0
; 
32'd20140: dataIn1 = 32'd1
; 
32'd20141: dataIn1 = 32'd2
; 
32'd20142: dataIn1 = 32'd5
; 
32'd20143: dataIn1 = 32'd11
; 
32'd20144: dataIn1 = 32'd13
; 
32'd20145: dataIn1 = 32'd17
; 
32'd20146: dataIn1 = 32'd19
; 
32'd20147: dataIn1 = 32'd20
; 
32'd20148: dataIn1 = 32'd23
; 
32'd20149: dataIn1 = 32'd25
; 
32'd20150: dataIn1 = 32'd28
; 
32'd20151: dataIn1 = 32'd30
; 
32'd20152: dataIn1 = 32'd34
; 
32'd20153: dataIn1 = 32'd35
; 
32'd20154: dataIn1 = 32'd36
; 
32'd20155: dataIn1 = 32'd39
; 
32'd20156: dataIn1 = 32'd40
; 
32'd20157: dataIn1 = 32'd42
; 
32'd20158: dataIn1 = 32'd43
; 
32'd20159: dataIn1 = 32'd56
; 
32'd20160: dataIn1 = 32'd62
; 
32'd20161: dataIn1 = 32'd63
; 
32'd20162: dataIn1 = 32'd1
; 
32'd20163: dataIn1 = 32'd2
; 
32'd20164: dataIn1 = 32'd7
; 
32'd20165: dataIn1 = 32'd9
; 
32'd20166: dataIn1 = 32'd11
; 
32'd20167: dataIn1 = 32'd18
; 
32'd20168: dataIn1 = 32'd19
; 
32'd20169: dataIn1 = 32'd22
; 
32'd20170: dataIn1 = 32'd28
; 
32'd20171: dataIn1 = 32'd30
; 
32'd20172: dataIn1 = 32'd32
; 
32'd20173: dataIn1 = 32'd34
; 
32'd20174: dataIn1 = 32'd35
; 
32'd20175: dataIn1 = 32'd36
; 
32'd20176: dataIn1 = 32'd38
; 
32'd20177: dataIn1 = 32'd39
; 
32'd20178: dataIn1 = 32'd43
; 
32'd20179: dataIn1 = 32'd50
; 
32'd20180: dataIn1 = 32'd56
; 
32'd20181: dataIn1 = 32'd61
; 
32'd20182: dataIn1 = 32'd5
; 
32'd20183: dataIn1 = 32'd6
; 
32'd20184: dataIn1 = 32'd9
; 
32'd20185: dataIn1 = 32'd10
; 
32'd20186: dataIn1 = 32'd12
; 
32'd20187: dataIn1 = 32'd15
; 
32'd20188: dataIn1 = 32'd17
; 
32'd20189: dataIn1 = 32'd27
; 
32'd20190: dataIn1 = 32'd32
; 
32'd20191: dataIn1 = 32'd33
; 
32'd20192: dataIn1 = 32'd34
; 
32'd20193: dataIn1 = 32'd35
; 
32'd20194: dataIn1 = 32'd39
; 
32'd20195: dataIn1 = 32'd40
; 
32'd20196: dataIn1 = 32'd41
; 
32'd20197: dataIn1 = 32'd42
; 
32'd20198: dataIn1 = 32'd43
; 
32'd20199: dataIn1 = 32'd45
; 
32'd20200: dataIn1 = 32'd47
; 
32'd20201: dataIn1 = 32'd48
; 
32'd20202: dataIn1 = 32'd49
; 
32'd20203: dataIn1 = 32'd50
; 
32'd20204: dataIn1 = 32'd54
; 
32'd20205: dataIn1 = 32'd55
; 
32'd20206: dataIn1 = 32'd60
; 
32'd20207: dataIn1 = 32'd63
; 
32'd20208: dataIn1 = 32'd1
; 
32'd20209: dataIn1 = 32'd2
; 
32'd20210: dataIn1 = 32'd10
; 
32'd20211: dataIn1 = 32'd11
; 
32'd20212: dataIn1 = 32'd12
; 
32'd20213: dataIn1 = 32'd14
; 
32'd20214: dataIn1 = 32'd18
; 
32'd20215: dataIn1 = 32'd22
; 
32'd20216: dataIn1 = 32'd23
; 
32'd20217: dataIn1 = 32'd28
; 
32'd20218: dataIn1 = 32'd29
; 
32'd20219: dataIn1 = 32'd30
; 
32'd20220: dataIn1 = 32'd34
; 
32'd20221: dataIn1 = 32'd41
; 
32'd20222: dataIn1 = 32'd42
; 
32'd20223: dataIn1 = 32'd43
; 
32'd20224: dataIn1 = 32'd44
; 
32'd20225: dataIn1 = 32'd49
; 
32'd20226: dataIn1 = 32'd52
; 
32'd20227: dataIn1 = 32'd53
; 
32'd20228: dataIn1 = 32'd54
; 
32'd20229: dataIn1 = 32'd56
; 
32'd20230: dataIn1 = 32'd58
; 
32'd20231: dataIn1 = 32'd61
; 
32'd20232: dataIn1 = 32'd0
; 
32'd20233: dataIn1 = 32'd2
; 
32'd20234: dataIn1 = 32'd5
; 
32'd20235: dataIn1 = 32'd6
; 
32'd20236: dataIn1 = 32'd11
; 
32'd20237: dataIn1 = 32'd14
; 
32'd20238: dataIn1 = 32'd15
; 
32'd20239: dataIn1 = 32'd18
; 
32'd20240: dataIn1 = 32'd19
; 
32'd20241: dataIn1 = 32'd22
; 
32'd20242: dataIn1 = 32'd26
; 
32'd20243: dataIn1 = 32'd31
; 
32'd20244: dataIn1 = 32'd32
; 
32'd20245: dataIn1 = 32'd35
; 
32'd20246: dataIn1 = 32'd36
; 
32'd20247: dataIn1 = 32'd41
; 
32'd20248: dataIn1 = 32'd47
; 
32'd20249: dataIn1 = 32'd48
; 
32'd20250: dataIn1 = 32'd50
; 
32'd20251: dataIn1 = 32'd53
; 
32'd20252: dataIn1 = 32'd54
; 
32'd20253: dataIn1 = 32'd58
; 
32'd20254: dataIn1 = 32'd62
; 
32'd20255: dataIn1 = 32'd63
; 
32'd20256: dataIn1 = 32'd1
; 
32'd20257: dataIn1 = 32'd2
; 
32'd20258: dataIn1 = 32'd3
; 
32'd20259: dataIn1 = 32'd4
; 
32'd20260: dataIn1 = 32'd7
; 
32'd20261: dataIn1 = 32'd13
; 
32'd20262: dataIn1 = 32'd14
; 
32'd20263: dataIn1 = 32'd15
; 
32'd20264: dataIn1 = 32'd20
; 
32'd20265: dataIn1 = 32'd22
; 
32'd20266: dataIn1 = 32'd24
; 
32'd20267: dataIn1 = 32'd25
; 
32'd20268: dataIn1 = 32'd29
; 
32'd20269: dataIn1 = 32'd32
; 
32'd20270: dataIn1 = 32'd34
; 
32'd20271: dataIn1 = 32'd36
; 
32'd20272: dataIn1 = 32'd38
; 
32'd20273: dataIn1 = 32'd39
; 
32'd20274: dataIn1 = 32'd42
; 
32'd20275: dataIn1 = 32'd43
; 
32'd20276: dataIn1 = 32'd47
; 
32'd20277: dataIn1 = 32'd49
; 
32'd20278: dataIn1 = 32'd50
; 
32'd20279: dataIn1 = 32'd53
; 
32'd20280: dataIn1 = 32'd54
; 
32'd20281: dataIn1 = 32'd60
; 
32'd20282: dataIn1 = 32'd0
; 
32'd20283: dataIn1 = 32'd6
; 
32'd20284: dataIn1 = 32'd7
; 
32'd20285: dataIn1 = 32'd14
; 
32'd20286: dataIn1 = 32'd16
; 
32'd20287: dataIn1 = 32'd18
; 
32'd20288: dataIn1 = 32'd19
; 
32'd20289: dataIn1 = 32'd21
; 
32'd20290: dataIn1 = 32'd24
; 
32'd20291: dataIn1 = 32'd25
; 
32'd20292: dataIn1 = 32'd28
; 
32'd20293: dataIn1 = 32'd30
; 
32'd20294: dataIn1 = 32'd32
; 
32'd20295: dataIn1 = 32'd33
; 
32'd20296: dataIn1 = 32'd34
; 
32'd20297: dataIn1 = 32'd35
; 
32'd20298: dataIn1 = 32'd39
; 
32'd20299: dataIn1 = 32'd43
; 
32'd20300: dataIn1 = 32'd47
; 
32'd20301: dataIn1 = 32'd48
; 
32'd20302: dataIn1 = 32'd51
; 
32'd20303: dataIn1 = 32'd53
; 
32'd20304: dataIn1 = 32'd56
; 
32'd20305: dataIn1 = 32'd59
; 
32'd20306: dataIn1 = 32'd60
; 
32'd20307: dataIn1 = 32'd62
; 
32'd20308: dataIn1 = 32'd63
; 
32'd20309: dataIn1 = 32'd2
; 
32'd20310: dataIn1 = 32'd6
; 
32'd20311: dataIn1 = 32'd7
; 
32'd20312: dataIn1 = 32'd9
; 
32'd20313: dataIn1 = 32'd11
; 
32'd20314: dataIn1 = 32'd13
; 
32'd20315: dataIn1 = 32'd14
; 
32'd20316: dataIn1 = 32'd15
; 
32'd20317: dataIn1 = 32'd20
; 
32'd20318: dataIn1 = 32'd22
; 
32'd20319: dataIn1 = 32'd26
; 
32'd20320: dataIn1 = 32'd27
; 
32'd20321: dataIn1 = 32'd33
; 
32'd20322: dataIn1 = 32'd36
; 
32'd20323: dataIn1 = 32'd38
; 
32'd20324: dataIn1 = 32'd40
; 
32'd20325: dataIn1 = 32'd44
; 
32'd20326: dataIn1 = 32'd46
; 
32'd20327: dataIn1 = 32'd47
; 
32'd20328: dataIn1 = 32'd48
; 
32'd20329: dataIn1 = 32'd49
; 
32'd20330: dataIn1 = 32'd51
; 
32'd20331: dataIn1 = 32'd52
; 
32'd20332: dataIn1 = 32'd56
; 
32'd20333: dataIn1 = 32'd57
; 
32'd20334: dataIn1 = 32'd58
; 
32'd20335: dataIn1 = 32'd3
; 
32'd20336: dataIn1 = 32'd5
; 
32'd20337: dataIn1 = 32'd9
; 
32'd20338: dataIn1 = 32'd13
; 
32'd20339: dataIn1 = 32'd16
; 
32'd20340: dataIn1 = 32'd21
; 
32'd20341: dataIn1 = 32'd23
; 
32'd20342: dataIn1 = 32'd25
; 
32'd20343: dataIn1 = 32'd28
; 
32'd20344: dataIn1 = 32'd31
; 
32'd20345: dataIn1 = 32'd33
; 
32'd20346: dataIn1 = 32'd35
; 
32'd20347: dataIn1 = 32'd38
; 
32'd20348: dataIn1 = 32'd43
; 
32'd20349: dataIn1 = 32'd44
; 
32'd20350: dataIn1 = 32'd50
; 
32'd20351: dataIn1 = 32'd52
; 
32'd20352: dataIn1 = 32'd53
; 
32'd20353: dataIn1 = 32'd56
; 
32'd20354: dataIn1 = 32'd60
; 
32'd20355: dataIn1 = 32'd61
; 
32'd20356: dataIn1 = 32'd62
; 
32'd20357: dataIn1 = 32'd63
; 
32'd20358: dataIn1 = 32'd1
; 
32'd20359: dataIn1 = 32'd2
; 
32'd20360: dataIn1 = 32'd5
; 
32'd20361: dataIn1 = 32'd6
; 
32'd20362: dataIn1 = 32'd7
; 
32'd20363: dataIn1 = 32'd8
; 
32'd20364: dataIn1 = 32'd9
; 
32'd20365: dataIn1 = 32'd14
; 
32'd20366: dataIn1 = 32'd16
; 
32'd20367: dataIn1 = 32'd19
; 
32'd20368: dataIn1 = 32'd20
; 
32'd20369: dataIn1 = 32'd21
; 
32'd20370: dataIn1 = 32'd27
; 
32'd20371: dataIn1 = 32'd30
; 
32'd20372: dataIn1 = 32'd31
; 
32'd20373: dataIn1 = 32'd33
; 
32'd20374: dataIn1 = 32'd34
; 
32'd20375: dataIn1 = 32'd36
; 
32'd20376: dataIn1 = 32'd39
; 
32'd20377: dataIn1 = 32'd40
; 
32'd20378: dataIn1 = 32'd41
; 
32'd20379: dataIn1 = 32'd44
; 
32'd20380: dataIn1 = 32'd52
; 
32'd20381: dataIn1 = 32'd57
; 
32'd20382: dataIn1 = 32'd62
; 
32'd20383: dataIn1 = 32'd63
; 
32'd20384: dataIn1 = 32'd5
; 
32'd20385: dataIn1 = 32'd9
; 
32'd20386: dataIn1 = 32'd10
; 
32'd20387: dataIn1 = 32'd19
; 
32'd20388: dataIn1 = 32'd20
; 
32'd20389: dataIn1 = 32'd21
; 
32'd20390: dataIn1 = 32'd22
; 
32'd20391: dataIn1 = 32'd26
; 
32'd20392: dataIn1 = 32'd30
; 
32'd20393: dataIn1 = 32'd31
; 
32'd20394: dataIn1 = 32'd32
; 
32'd20395: dataIn1 = 32'd34
; 
32'd20396: dataIn1 = 32'd38
; 
32'd20397: dataIn1 = 32'd39
; 
32'd20398: dataIn1 = 32'd41
; 
32'd20399: dataIn1 = 32'd42
; 
32'd20400: dataIn1 = 32'd45
; 
32'd20401: dataIn1 = 32'd46
; 
32'd20402: dataIn1 = 32'd50
; 
32'd20403: dataIn1 = 32'd51
; 
32'd20404: dataIn1 = 32'd52
; 
32'd20405: dataIn1 = 32'd53
; 
32'd20406: dataIn1 = 32'd54
; 
32'd20407: dataIn1 = 32'd59
; 
32'd20408: dataIn1 = 32'd61
; 
32'd20409: dataIn1 = 32'd0
; 
32'd20410: dataIn1 = 32'd1
; 
32'd20411: dataIn1 = 32'd8
; 
32'd20412: dataIn1 = 32'd17
; 
32'd20413: dataIn1 = 32'd18
; 
32'd20414: dataIn1 = 32'd20
; 
32'd20415: dataIn1 = 32'd24
; 
32'd20416: dataIn1 = 32'd27
; 
32'd20417: dataIn1 = 32'd32
; 
32'd20418: dataIn1 = 32'd38
; 
32'd20419: dataIn1 = 32'd39
; 
32'd20420: dataIn1 = 32'd41
; 
32'd20421: dataIn1 = 32'd42
; 
32'd20422: dataIn1 = 32'd44
; 
32'd20423: dataIn1 = 32'd48
; 
32'd20424: dataIn1 = 32'd56
; 
32'd20425: dataIn1 = 32'd57
; 
32'd20426: dataIn1 = 32'd60
; 
32'd20427: dataIn1 = 32'd0
; 
32'd20428: dataIn1 = 32'd1
; 
32'd20429: dataIn1 = 32'd3
; 
32'd20430: dataIn1 = 32'd8
; 
32'd20431: dataIn1 = 32'd9
; 
32'd20432: dataIn1 = 32'd11
; 
32'd20433: dataIn1 = 32'd12
; 
32'd20434: dataIn1 = 32'd20
; 
32'd20435: dataIn1 = 32'd21
; 
32'd20436: dataIn1 = 32'd28
; 
32'd20437: dataIn1 = 32'd29
; 
32'd20438: dataIn1 = 32'd32
; 
32'd20439: dataIn1 = 32'd34
; 
32'd20440: dataIn1 = 32'd35
; 
32'd20441: dataIn1 = 32'd39
; 
32'd20442: dataIn1 = 32'd44
; 
32'd20443: dataIn1 = 32'd45
; 
32'd20444: dataIn1 = 32'd51
; 
32'd20445: dataIn1 = 32'd52
; 
32'd20446: dataIn1 = 32'd53
; 
32'd20447: dataIn1 = 32'd55
; 
32'd20448: dataIn1 = 32'd56
; 
32'd20449: dataIn1 = 32'd61
; 
32'd20450: dataIn1 = 32'd62
; 
32'd20451: dataIn1 = 32'd0
; 
32'd20452: dataIn1 = 32'd7
; 
32'd20453: dataIn1 = 32'd11
; 
32'd20454: dataIn1 = 32'd21
; 
32'd20455: dataIn1 = 32'd25
; 
32'd20456: dataIn1 = 32'd26
; 
32'd20457: dataIn1 = 32'd36
; 
32'd20458: dataIn1 = 32'd38
; 
32'd20459: dataIn1 = 32'd39
; 
32'd20460: dataIn1 = 32'd42
; 
32'd20461: dataIn1 = 32'd44
; 
32'd20462: dataIn1 = 32'd48
; 
32'd20463: dataIn1 = 32'd49
; 
32'd20464: dataIn1 = 32'd50
; 
32'd20465: dataIn1 = 32'd52
; 
32'd20466: dataIn1 = 32'd53
; 
32'd20467: dataIn1 = 32'd54
; 
32'd20468: dataIn1 = 32'd55
; 
32'd20469: dataIn1 = 32'd58
; 
32'd20470: dataIn1 = 32'd61
; 
32'd20471: dataIn1 = 32'd1
; 
32'd20472: dataIn1 = 32'd2
; 
32'd20473: dataIn1 = 32'd7
; 
32'd20474: dataIn1 = 32'd8
; 
32'd20475: dataIn1 = 32'd11
; 
32'd20476: dataIn1 = 32'd12
; 
32'd20477: dataIn1 = 32'd19
; 
32'd20478: dataIn1 = 32'd22
; 
32'd20479: dataIn1 = 32'd27
; 
32'd20480: dataIn1 = 32'd33
; 
32'd20481: dataIn1 = 32'd34
; 
32'd20482: dataIn1 = 32'd38
; 
32'd20483: dataIn1 = 32'd41
; 
32'd20484: dataIn1 = 32'd43
; 
32'd20485: dataIn1 = 32'd44
; 
32'd20486: dataIn1 = 32'd45
; 
32'd20487: dataIn1 = 32'd47
; 
32'd20488: dataIn1 = 32'd49
; 
32'd20489: dataIn1 = 32'd51
; 
32'd20490: dataIn1 = 32'd52
; 
32'd20491: dataIn1 = 32'd54
; 
32'd20492: dataIn1 = 32'd55
; 
32'd20493: dataIn1 = 32'd60
; 
32'd20494: dataIn1 = 32'd62
; 
32'd20495: dataIn1 = 32'd0
; 
32'd20496: dataIn1 = 32'd1
; 
32'd20497: dataIn1 = 32'd2
; 
32'd20498: dataIn1 = 32'd3
; 
32'd20499: dataIn1 = 32'd5
; 
32'd20500: dataIn1 = 32'd8
; 
32'd20501: dataIn1 = 32'd9
; 
32'd20502: dataIn1 = 32'd10
; 
32'd20503: dataIn1 = 32'd17
; 
32'd20504: dataIn1 = 32'd19
; 
32'd20505: dataIn1 = 32'd20
; 
32'd20506: dataIn1 = 32'd22
; 
32'd20507: dataIn1 = 32'd23
; 
32'd20508: dataIn1 = 32'd25
; 
32'd20509: dataIn1 = 32'd26
; 
32'd20510: dataIn1 = 32'd28
; 
32'd20511: dataIn1 = 32'd30
; 
32'd20512: dataIn1 = 32'd32
; 
32'd20513: dataIn1 = 32'd36
; 
32'd20514: dataIn1 = 32'd46
; 
32'd20515: dataIn1 = 32'd51
; 
32'd20516: dataIn1 = 32'd56
; 
32'd20517: dataIn1 = 32'd58
; 
32'd20518: dataIn1 = 32'd59
; 
32'd20519: dataIn1 = 32'd1
; 
32'd20520: dataIn1 = 32'd3
; 
32'd20521: dataIn1 = 32'd5
; 
32'd20522: dataIn1 = 32'd7
; 
32'd20523: dataIn1 = 32'd15
; 
32'd20524: dataIn1 = 32'd17
; 
32'd20525: dataIn1 = 32'd21
; 
32'd20526: dataIn1 = 32'd23
; 
32'd20527: dataIn1 = 32'd28
; 
32'd20528: dataIn1 = 32'd29
; 
32'd20529: dataIn1 = 32'd38
; 
32'd20530: dataIn1 = 32'd39
; 
32'd20531: dataIn1 = 32'd40
; 
32'd20532: dataIn1 = 32'd42
; 
32'd20533: dataIn1 = 32'd45
; 
32'd20534: dataIn1 = 32'd47
; 
32'd20535: dataIn1 = 32'd49
; 
32'd20536: dataIn1 = 32'd52
; 
32'd20537: dataIn1 = 32'd53
; 
32'd20538: dataIn1 = 32'd56
; 
32'd20539: dataIn1 = 32'd59
; 
32'd20540: dataIn1 = 32'd60
; 
32'd20541: dataIn1 = 32'd63
; 
32'd20542: dataIn1 = 32'd2
; 
32'd20543: dataIn1 = 32'd4
; 
32'd20544: dataIn1 = 32'd5
; 
32'd20545: dataIn1 = 32'd6
; 
32'd20546: dataIn1 = 32'd7
; 
32'd20547: dataIn1 = 32'd9
; 
32'd20548: dataIn1 = 32'd10
; 
32'd20549: dataIn1 = 32'd11
; 
32'd20550: dataIn1 = 32'd15
; 
32'd20551: dataIn1 = 32'd19
; 
32'd20552: dataIn1 = 32'd23
; 
32'd20553: dataIn1 = 32'd24
; 
32'd20554: dataIn1 = 32'd25
; 
32'd20555: dataIn1 = 32'd26
; 
32'd20556: dataIn1 = 32'd27
; 
32'd20557: dataIn1 = 32'd31
; 
32'd20558: dataIn1 = 32'd33
; 
32'd20559: dataIn1 = 32'd34
; 
32'd20560: dataIn1 = 32'd37
; 
32'd20561: dataIn1 = 32'd41
; 
32'd20562: dataIn1 = 32'd42
; 
32'd20563: dataIn1 = 32'd44
; 
32'd20564: dataIn1 = 32'd45
; 
32'd20565: dataIn1 = 32'd47
; 
32'd20566: dataIn1 = 32'd51
; 
32'd20567: dataIn1 = 32'd52
; 
32'd20568: dataIn1 = 32'd55
; 
32'd20569: dataIn1 = 32'd56
; 
32'd20570: dataIn1 = 32'd61
; 
32'd20571: dataIn1 = 32'd63
; 
32'd20572: dataIn1 = 32'd2
; 
32'd20573: dataIn1 = 32'd4
; 
32'd20574: dataIn1 = 32'd5
; 
32'd20575: dataIn1 = 32'd8
; 
32'd20576: dataIn1 = 32'd9
; 
32'd20577: dataIn1 = 32'd14
; 
32'd20578: dataIn1 = 32'd19
; 
32'd20579: dataIn1 = 32'd20
; 
32'd20580: dataIn1 = 32'd21
; 
32'd20581: dataIn1 = 32'd22
; 
32'd20582: dataIn1 = 32'd23
; 
32'd20583: dataIn1 = 32'd24
; 
32'd20584: dataIn1 = 32'd26
; 
32'd20585: dataIn1 = 32'd27
; 
32'd20586: dataIn1 = 32'd29
; 
32'd20587: dataIn1 = 32'd32
; 
32'd20588: dataIn1 = 32'd33
; 
32'd20589: dataIn1 = 32'd35
; 
32'd20590: dataIn1 = 32'd40
; 
32'd20591: dataIn1 = 32'd42
; 
32'd20592: dataIn1 = 32'd46
; 
32'd20593: dataIn1 = 32'd48
; 
32'd20594: dataIn1 = 32'd49
; 
32'd20595: dataIn1 = 32'd51
; 
32'd20596: dataIn1 = 32'd52
; 
32'd20597: dataIn1 = 32'd56
; 
32'd20598: dataIn1 = 32'd57
; 
32'd20599: dataIn1 = 32'd58
; 
32'd20600: dataIn1 = 32'd60
; 
32'd20601: dataIn1 = 32'd2
; 
32'd20602: dataIn1 = 32'd7
; 
32'd20603: dataIn1 = 32'd8
; 
32'd20604: dataIn1 = 32'd9
; 
32'd20605: dataIn1 = 32'd12
; 
32'd20606: dataIn1 = 32'd13
; 
32'd20607: dataIn1 = 32'd15
; 
32'd20608: dataIn1 = 32'd16
; 
32'd20609: dataIn1 = 32'd25
; 
32'd20610: dataIn1 = 32'd26
; 
32'd20611: dataIn1 = 32'd35
; 
32'd20612: dataIn1 = 32'd37
; 
32'd20613: dataIn1 = 32'd38
; 
32'd20614: dataIn1 = 32'd39
; 
32'd20615: dataIn1 = 32'd42
; 
32'd20616: dataIn1 = 32'd48
; 
32'd20617: dataIn1 = 32'd49
; 
32'd20618: dataIn1 = 32'd50
; 
32'd20619: dataIn1 = 32'd51
; 
32'd20620: dataIn1 = 32'd53
; 
32'd20621: dataIn1 = 32'd58
; 
32'd20622: dataIn1 = 32'd60
; 
32'd20623: dataIn1 = 32'd0
; 
32'd20624: dataIn1 = 32'd2
; 
32'd20625: dataIn1 = 32'd3
; 
32'd20626: dataIn1 = 32'd5
; 
32'd20627: dataIn1 = 32'd8
; 
32'd20628: dataIn1 = 32'd9
; 
32'd20629: dataIn1 = 32'd10
; 
32'd20630: dataIn1 = 32'd11
; 
32'd20631: dataIn1 = 32'd12
; 
32'd20632: dataIn1 = 32'd14
; 
32'd20633: dataIn1 = 32'd18
; 
32'd20634: dataIn1 = 32'd19
; 
32'd20635: dataIn1 = 32'd21
; 
32'd20636: dataIn1 = 32'd23
; 
32'd20637: dataIn1 = 32'd25
; 
32'd20638: dataIn1 = 32'd27
; 
32'd20639: dataIn1 = 32'd31
; 
32'd20640: dataIn1 = 32'd36
; 
32'd20641: dataIn1 = 32'd44
; 
32'd20642: dataIn1 = 32'd49
; 
32'd20643: dataIn1 = 32'd54
; 
32'd20644: dataIn1 = 32'd57
; 
32'd20645: dataIn1 = 32'd60
; 
32'd20646: dataIn1 = 32'd1
; 
32'd20647: dataIn1 = 32'd8
; 
32'd20648: dataIn1 = 32'd11
; 
32'd20649: dataIn1 = 32'd12
; 
32'd20650: dataIn1 = 32'd16
; 
32'd20651: dataIn1 = 32'd18
; 
32'd20652: dataIn1 = 32'd21
; 
32'd20653: dataIn1 = 32'd22
; 
32'd20654: dataIn1 = 32'd24
; 
32'd20655: dataIn1 = 32'd27
; 
32'd20656: dataIn1 = 32'd34
; 
32'd20657: dataIn1 = 32'd36
; 
32'd20658: dataIn1 = 32'd37
; 
32'd20659: dataIn1 = 32'd44
; 
32'd20660: dataIn1 = 32'd45
; 
32'd20661: dataIn1 = 32'd50
; 
32'd20662: dataIn1 = 32'd51
; 
32'd20663: dataIn1 = 32'd54
; 
32'd20664: dataIn1 = 32'd58
; 
32'd20665: dataIn1 = 32'd0
; 
32'd20666: dataIn1 = 32'd1
; 
32'd20667: dataIn1 = 32'd3
; 
32'd20668: dataIn1 = 32'd4
; 
32'd20669: dataIn1 = 32'd6
; 
32'd20670: dataIn1 = 32'd12
; 
32'd20671: dataIn1 = 32'd14
; 
32'd20672: dataIn1 = 32'd15
; 
32'd20673: dataIn1 = 32'd18
; 
32'd20674: dataIn1 = 32'd21
; 
32'd20675: dataIn1 = 32'd25
; 
32'd20676: dataIn1 = 32'd26
; 
32'd20677: dataIn1 = 32'd27
; 
32'd20678: dataIn1 = 32'd28
; 
32'd20679: dataIn1 = 32'd29
; 
32'd20680: dataIn1 = 32'd32
; 
32'd20681: dataIn1 = 32'd40
; 
32'd20682: dataIn1 = 32'd42
; 
32'd20683: dataIn1 = 32'd44
; 
32'd20684: dataIn1 = 32'd47
; 
32'd20685: dataIn1 = 32'd50
; 
32'd20686: dataIn1 = 32'd52
; 
32'd20687: dataIn1 = 32'd54
; 
32'd20688: dataIn1 = 32'd57
; 
32'd20689: dataIn1 = 32'd61
; 
32'd20690: dataIn1 = 32'd62
; 
32'd20691: dataIn1 = 32'd63
; 
32'd20692: dataIn1 = 32'd3
; 
32'd20693: dataIn1 = 32'd4
; 
32'd20694: dataIn1 = 32'd5
; 
32'd20695: dataIn1 = 32'd12
; 
32'd20696: dataIn1 = 32'd22
; 
32'd20697: dataIn1 = 32'd26
; 
32'd20698: dataIn1 = 32'd28
; 
32'd20699: dataIn1 = 32'd30
; 
32'd20700: dataIn1 = 32'd32
; 
32'd20701: dataIn1 = 32'd33
; 
32'd20702: dataIn1 = 32'd34
; 
32'd20703: dataIn1 = 32'd35
; 
32'd20704: dataIn1 = 32'd38
; 
32'd20705: dataIn1 = 32'd40
; 
32'd20706: dataIn1 = 32'd41
; 
32'd20707: dataIn1 = 32'd43
; 
32'd20708: dataIn1 = 32'd44
; 
32'd20709: dataIn1 = 32'd47
; 
32'd20710: dataIn1 = 32'd52
; 
32'd20711: dataIn1 = 32'd53
; 
32'd20712: dataIn1 = 32'd54
; 
32'd20713: dataIn1 = 32'd56
; 
32'd20714: dataIn1 = 32'd59
; 
32'd20715: dataIn1 = 32'd60
; 
32'd20716: dataIn1 = 32'd61
; 
32'd20717: dataIn1 = 32'd3
; 
32'd20718: dataIn1 = 32'd6
; 
32'd20719: dataIn1 = 32'd9
; 
32'd20720: dataIn1 = 32'd10
; 
32'd20721: dataIn1 = 32'd12
; 
32'd20722: dataIn1 = 32'd13
; 
32'd20723: dataIn1 = 32'd14
; 
32'd20724: dataIn1 = 32'd15
; 
32'd20725: dataIn1 = 32'd17
; 
32'd20726: dataIn1 = 32'd21
; 
32'd20727: dataIn1 = 32'd22
; 
32'd20728: dataIn1 = 32'd25
; 
32'd20729: dataIn1 = 32'd26
; 
32'd20730: dataIn1 = 32'd28
; 
32'd20731: dataIn1 = 32'd31
; 
32'd20732: dataIn1 = 32'd36
; 
32'd20733: dataIn1 = 32'd38
; 
32'd20734: dataIn1 = 32'd43
; 
32'd20735: dataIn1 = 32'd52
; 
32'd20736: dataIn1 = 32'd55
; 
32'd20737: dataIn1 = 32'd57
; 
32'd20738: dataIn1 = 32'd60
; 
32'd20739: dataIn1 = 32'd62
; 
32'd20740: dataIn1 = 32'd0
; 
32'd20741: dataIn1 = 32'd1
; 
32'd20742: dataIn1 = 32'd4
; 
32'd20743: dataIn1 = 32'd5
; 
32'd20744: dataIn1 = 32'd9
; 
32'd20745: dataIn1 = 32'd14
; 
32'd20746: dataIn1 = 32'd19
; 
32'd20747: dataIn1 = 32'd23
; 
32'd20748: dataIn1 = 32'd30
; 
32'd20749: dataIn1 = 32'd31
; 
32'd20750: dataIn1 = 32'd33
; 
32'd20751: dataIn1 = 32'd38
; 
32'd20752: dataIn1 = 32'd39
; 
32'd20753: dataIn1 = 32'd42
; 
32'd20754: dataIn1 = 32'd43
; 
32'd20755: dataIn1 = 32'd46
; 
32'd20756: dataIn1 = 32'd51
; 
32'd20757: dataIn1 = 32'd55
; 
32'd20758: dataIn1 = 32'd62
; 
32'd20759: dataIn1 = 32'd2
; 
32'd20760: dataIn1 = 32'd4
; 
32'd20761: dataIn1 = 32'd5
; 
32'd20762: dataIn1 = 32'd14
; 
32'd20763: dataIn1 = 32'd17
; 
32'd20764: dataIn1 = 32'd20
; 
32'd20765: dataIn1 = 32'd21
; 
32'd20766: dataIn1 = 32'd23
; 
32'd20767: dataIn1 = 32'd25
; 
32'd20768: dataIn1 = 32'd26
; 
32'd20769: dataIn1 = 32'd33
; 
32'd20770: dataIn1 = 32'd36
; 
32'd20771: dataIn1 = 32'd49
; 
32'd20772: dataIn1 = 32'd52
; 
32'd20773: dataIn1 = 32'd57
; 
32'd20774: dataIn1 = 32'd59
; 
32'd20775: dataIn1 = 32'd60
; 
32'd20776: dataIn1 = 32'd62
; 
32'd20777: dataIn1 = 32'd1
; 
32'd20778: dataIn1 = 32'd3
; 
32'd20779: dataIn1 = 32'd11
; 
32'd20780: dataIn1 = 32'd18
; 
32'd20781: dataIn1 = 32'd22
; 
32'd20782: dataIn1 = 32'd24
; 
32'd20783: dataIn1 = 32'd26
; 
32'd20784: dataIn1 = 32'd30
; 
32'd20785: dataIn1 = 32'd32
; 
32'd20786: dataIn1 = 32'd33
; 
32'd20787: dataIn1 = 32'd36
; 
32'd20788: dataIn1 = 32'd37
; 
32'd20789: dataIn1 = 32'd38
; 
32'd20790: dataIn1 = 32'd39
; 
32'd20791: dataIn1 = 32'd40
; 
32'd20792: dataIn1 = 32'd42
; 
32'd20793: dataIn1 = 32'd48
; 
32'd20794: dataIn1 = 32'd50
; 
32'd20795: dataIn1 = 32'd53
; 
32'd20796: dataIn1 = 32'd55
; 
32'd20797: dataIn1 = 32'd57
; 
32'd20798: dataIn1 = 32'd58
; 
32'd20799: dataIn1 = 32'd62
; 
32'd20800: dataIn1 = 32'd63
; 
32'd20801: dataIn1 = 32'd1
; 
32'd20802: dataIn1 = 32'd7
; 
32'd20803: dataIn1 = 32'd8
; 
32'd20804: dataIn1 = 32'd9
; 
32'd20805: dataIn1 = 32'd11
; 
32'd20806: dataIn1 = 32'd13
; 
32'd20807: dataIn1 = 32'd15
; 
32'd20808: dataIn1 = 32'd21
; 
32'd20809: dataIn1 = 32'd22
; 
32'd20810: dataIn1 = 32'd23
; 
32'd20811: dataIn1 = 32'd24
; 
32'd20812: dataIn1 = 32'd29
; 
32'd20813: dataIn1 = 32'd32
; 
32'd20814: dataIn1 = 32'd36
; 
32'd20815: dataIn1 = 32'd38
; 
32'd20816: dataIn1 = 32'd41
; 
32'd20817: dataIn1 = 32'd42
; 
32'd20818: dataIn1 = 32'd50
; 
32'd20819: dataIn1 = 32'd53
; 
32'd20820: dataIn1 = 32'd55
; 
32'd20821: dataIn1 = 32'd56
; 
32'd20822: dataIn1 = 32'd58
; 
32'd20823: dataIn1 = 32'd60
; 
32'd20824: dataIn1 = 32'd61
; 
32'd20825: dataIn1 = 32'd2
; 
32'd20826: dataIn1 = 32'd3
; 
32'd20827: dataIn1 = 32'd4
; 
32'd20828: dataIn1 = 32'd8
; 
32'd20829: dataIn1 = 32'd11
; 
32'd20830: dataIn1 = 32'd16
; 
32'd20831: dataIn1 = 32'd17
; 
32'd20832: dataIn1 = 32'd18
; 
32'd20833: dataIn1 = 32'd19
; 
32'd20834: dataIn1 = 32'd24
; 
32'd20835: dataIn1 = 32'd25
; 
32'd20836: dataIn1 = 32'd28
; 
32'd20837: dataIn1 = 32'd30
; 
32'd20838: dataIn1 = 32'd32
; 
32'd20839: dataIn1 = 32'd35
; 
32'd20840: dataIn1 = 32'd36
; 
32'd20841: dataIn1 = 32'd39
; 
32'd20842: dataIn1 = 32'd41
; 
32'd20843: dataIn1 = 32'd44
; 
32'd20844: dataIn1 = 32'd46
; 
32'd20845: dataIn1 = 32'd48
; 
32'd20846: dataIn1 = 32'd51
; 
32'd20847: dataIn1 = 32'd57
; 
32'd20848: dataIn1 = 32'd58
; 
32'd20849: dataIn1 = 32'd59
; 
32'd20850: dataIn1 = 32'd63
; 
32'd20851: dataIn1 = 32'd0
; 
32'd20852: dataIn1 = 32'd5
; 
32'd20853: dataIn1 = 32'd6
; 
32'd20854: dataIn1 = 32'd11
; 
32'd20855: dataIn1 = 32'd12
; 
32'd20856: dataIn1 = 32'd13
; 
32'd20857: dataIn1 = 32'd14
; 
32'd20858: dataIn1 = 32'd15
; 
32'd20859: dataIn1 = 32'd20
; 
32'd20860: dataIn1 = 32'd21
; 
32'd20861: dataIn1 = 32'd24
; 
32'd20862: dataIn1 = 32'd26
; 
32'd20863: dataIn1 = 32'd35
; 
32'd20864: dataIn1 = 32'd36
; 
32'd20865: dataIn1 = 32'd38
; 
32'd20866: dataIn1 = 32'd44
; 
32'd20867: dataIn1 = 32'd45
; 
32'd20868: dataIn1 = 32'd46
; 
32'd20869: dataIn1 = 32'd47
; 
32'd20870: dataIn1 = 32'd48
; 
32'd20871: dataIn1 = 32'd50
; 
32'd20872: dataIn1 = 32'd54
; 
32'd20873: dataIn1 = 32'd55
; 
32'd20874: dataIn1 = 32'd57
; 
32'd20875: dataIn1 = 32'd62
; 
32'd20876: dataIn1 = 32'd0
; 
32'd20877: dataIn1 = 32'd1
; 
32'd20878: dataIn1 = 32'd4
; 
32'd20879: dataIn1 = 32'd7
; 
32'd20880: dataIn1 = 32'd8
; 
32'd20881: dataIn1 = 32'd12
; 
32'd20882: dataIn1 = 32'd14
; 
32'd20883: dataIn1 = 32'd21
; 
32'd20884: dataIn1 = 32'd22
; 
32'd20885: dataIn1 = 32'd23
; 
32'd20886: dataIn1 = 32'd24
; 
32'd20887: dataIn1 = 32'd28
; 
32'd20888: dataIn1 = 32'd29
; 
32'd20889: dataIn1 = 32'd33
; 
32'd20890: dataIn1 = 32'd37
; 
32'd20891: dataIn1 = 32'd40
; 
32'd20892: dataIn1 = 32'd41
; 
32'd20893: dataIn1 = 32'd49
; 
32'd20894: dataIn1 = 32'd56
; 
32'd20895: dataIn1 = 32'd58
; 
32'd20896: dataIn1 = 32'd60
; 
32'd20897: dataIn1 = 32'd1
; 
32'd20898: dataIn1 = 32'd3
; 
32'd20899: dataIn1 = 32'd7
; 
32'd20900: dataIn1 = 32'd8
; 
32'd20901: dataIn1 = 32'd11
; 
32'd20902: dataIn1 = 32'd14
; 
32'd20903: dataIn1 = 32'd16
; 
32'd20904: dataIn1 = 32'd18
; 
32'd20905: dataIn1 = 32'd23
; 
32'd20906: dataIn1 = 32'd25
; 
32'd20907: dataIn1 = 32'd26
; 
32'd20908: dataIn1 = 32'd31
; 
32'd20909: dataIn1 = 32'd32
; 
32'd20910: dataIn1 = 32'd34
; 
32'd20911: dataIn1 = 32'd37
; 
32'd20912: dataIn1 = 32'd39
; 
32'd20913: dataIn1 = 32'd40
; 
32'd20914: dataIn1 = 32'd47
; 
32'd20915: dataIn1 = 32'd49
; 
32'd20916: dataIn1 = 32'd50
; 
32'd20917: dataIn1 = 32'd52
; 
32'd20918: dataIn1 = 32'd54
; 
32'd20919: dataIn1 = 32'd56
; 
32'd20920: dataIn1 = 32'd63
; 
32'd20921: dataIn1 = 32'd2
; 
32'd20922: dataIn1 = 32'd4
; 
32'd20923: dataIn1 = 32'd15
; 
32'd20924: dataIn1 = 32'd16
; 
32'd20925: dataIn1 = 32'd18
; 
32'd20926: dataIn1 = 32'd25
; 
32'd20927: dataIn1 = 32'd26
; 
32'd20928: dataIn1 = 32'd27
; 
32'd20929: dataIn1 = 32'd32
; 
32'd20930: dataIn1 = 32'd34
; 
32'd20931: dataIn1 = 32'd36
; 
32'd20932: dataIn1 = 32'd37
; 
32'd20933: dataIn1 = 32'd39
; 
32'd20934: dataIn1 = 32'd42
; 
32'd20935: dataIn1 = 32'd51
; 
32'd20936: dataIn1 = 32'd57
; 
32'd20937: dataIn1 = 32'd60
; 
32'd20938: dataIn1 = 32'd63
; 
32'd20939: dataIn1 = 32'd0
; 
32'd20940: dataIn1 = 32'd2
; 
32'd20941: dataIn1 = 32'd3
; 
32'd20942: dataIn1 = 32'd5
; 
32'd20943: dataIn1 = 32'd6
; 
32'd20944: dataIn1 = 32'd8
; 
32'd20945: dataIn1 = 32'd11
; 
32'd20946: dataIn1 = 32'd13
; 
32'd20947: dataIn1 = 32'd16
; 
32'd20948: dataIn1 = 32'd18
; 
32'd20949: dataIn1 = 32'd22
; 
32'd20950: dataIn1 = 32'd32
; 
32'd20951: dataIn1 = 32'd33
; 
32'd20952: dataIn1 = 32'd44
; 
32'd20953: dataIn1 = 32'd45
; 
32'd20954: dataIn1 = 32'd50
; 
32'd20955: dataIn1 = 32'd51
; 
32'd20956: dataIn1 = 32'd52
; 
32'd20957: dataIn1 = 32'd58
; 
32'd20958: dataIn1 = 32'd62
; 
32'd20959: dataIn1 = 32'd63
; 
32'd20960: dataIn1 = 32'd0
; 
32'd20961: dataIn1 = 32'd3
; 
32'd20962: dataIn1 = 32'd7
; 
32'd20963: dataIn1 = 32'd12
; 
32'd20964: dataIn1 = 32'd14
; 
32'd20965: dataIn1 = 32'd17
; 
32'd20966: dataIn1 = 32'd19
; 
32'd20967: dataIn1 = 32'd20
; 
32'd20968: dataIn1 = 32'd22
; 
32'd20969: dataIn1 = 32'd27
; 
32'd20970: dataIn1 = 32'd30
; 
32'd20971: dataIn1 = 32'd36
; 
32'd20972: dataIn1 = 32'd37
; 
32'd20973: dataIn1 = 32'd38
; 
32'd20974: dataIn1 = 32'd49
; 
32'd20975: dataIn1 = 32'd51
; 
32'd20976: dataIn1 = 32'd53
; 
32'd20977: dataIn1 = 32'd54
; 
32'd20978: dataIn1 = 32'd55
; 
32'd20979: dataIn1 = 32'd58
; 
32'd20980: dataIn1 = 32'd61
; 
32'd20981: dataIn1 = 32'd1
; 
32'd20982: dataIn1 = 32'd2
; 
32'd20983: dataIn1 = 32'd6
; 
32'd20984: dataIn1 = 32'd7
; 
32'd20985: dataIn1 = 32'd9
; 
32'd20986: dataIn1 = 32'd11
; 
32'd20987: dataIn1 = 32'd12
; 
32'd20988: dataIn1 = 32'd13
; 
32'd20989: dataIn1 = 32'd14
; 
32'd20990: dataIn1 = 32'd15
; 
32'd20991: dataIn1 = 32'd17
; 
32'd20992: dataIn1 = 32'd18
; 
32'd20993: dataIn1 = 32'd20
; 
32'd20994: dataIn1 = 32'd21
; 
32'd20995: dataIn1 = 32'd22
; 
32'd20996: dataIn1 = 32'd23
; 
32'd20997: dataIn1 = 32'd24
; 
32'd20998: dataIn1 = 32'd28
; 
32'd20999: dataIn1 = 32'd29
; 
32'd21000: dataIn1 = 32'd32
; 
32'd21001: dataIn1 = 32'd38
; 
32'd21002: dataIn1 = 32'd39
; 
32'd21003: dataIn1 = 32'd40
; 
32'd21004: dataIn1 = 32'd42
; 
32'd21005: dataIn1 = 32'd47
; 
32'd21006: dataIn1 = 32'd55
; 
32'd21007: dataIn1 = 32'd58
; 
32'd21008: dataIn1 = 32'd61
; 
32'd21009: dataIn1 = 32'd62
; 
32'd21010: dataIn1 = 32'd0
; 
32'd21011: dataIn1 = 32'd1
; 
32'd21012: dataIn1 = 32'd3
; 
32'd21013: dataIn1 = 32'd5
; 
32'd21014: dataIn1 = 32'd6
; 
32'd21015: dataIn1 = 32'd8
; 
32'd21016: dataIn1 = 32'd10
; 
32'd21017: dataIn1 = 32'd11
; 
32'd21018: dataIn1 = 32'd15
; 
32'd21019: dataIn1 = 32'd16
; 
32'd21020: dataIn1 = 32'd21
; 
32'd21021: dataIn1 = 32'd23
; 
32'd21022: dataIn1 = 32'd25
; 
32'd21023: dataIn1 = 32'd27
; 
32'd21024: dataIn1 = 32'd35
; 
32'd21025: dataIn1 = 32'd36
; 
32'd21026: dataIn1 = 32'd38
; 
32'd21027: dataIn1 = 32'd41
; 
32'd21028: dataIn1 = 32'd42
; 
32'd21029: dataIn1 = 32'd43
; 
32'd21030: dataIn1 = 32'd48
; 
32'd21031: dataIn1 = 32'd51
; 
32'd21032: dataIn1 = 32'd53
; 
32'd21033: dataIn1 = 32'd55
; 
32'd21034: dataIn1 = 32'd56
; 
32'd21035: dataIn1 = 32'd58
; 
32'd21036: dataIn1 = 32'd61
; 
32'd21037: dataIn1 = 32'd63
; 
32'd21038: dataIn1 = 32'd1
; 
32'd21039: dataIn1 = 32'd2
; 
32'd21040: dataIn1 = 32'd3
; 
32'd21041: dataIn1 = 32'd5
; 
32'd21042: dataIn1 = 32'd8
; 
32'd21043: dataIn1 = 32'd10
; 
32'd21044: dataIn1 = 32'd11
; 
32'd21045: dataIn1 = 32'd12
; 
32'd21046: dataIn1 = 32'd14
; 
32'd21047: dataIn1 = 32'd15
; 
32'd21048: dataIn1 = 32'd19
; 
32'd21049: dataIn1 = 32'd22
; 
32'd21050: dataIn1 = 32'd24
; 
32'd21051: dataIn1 = 32'd28
; 
32'd21052: dataIn1 = 32'd30
; 
32'd21053: dataIn1 = 32'd31
; 
32'd21054: dataIn1 = 32'd32
; 
32'd21055: dataIn1 = 32'd33
; 
32'd21056: dataIn1 = 32'd41
; 
32'd21057: dataIn1 = 32'd43
; 
32'd21058: dataIn1 = 32'd45
; 
32'd21059: dataIn1 = 32'd47
; 
32'd21060: dataIn1 = 32'd48
; 
32'd21061: dataIn1 = 32'd49
; 
32'd21062: dataIn1 = 32'd51
; 
32'd21063: dataIn1 = 32'd53
; 
32'd21064: dataIn1 = 32'd57
; 
32'd21065: dataIn1 = 32'd58
; 
32'd21066: dataIn1 = 32'd62
; 
32'd21067: dataIn1 = 32'd0
; 
32'd21068: dataIn1 = 32'd3
; 
32'd21069: dataIn1 = 32'd12
; 
32'd21070: dataIn1 = 32'd15
; 
32'd21071: dataIn1 = 32'd16
; 
32'd21072: dataIn1 = 32'd22
; 
32'd21073: dataIn1 = 32'd25
; 
32'd21074: dataIn1 = 32'd27
; 
32'd21075: dataIn1 = 32'd29
; 
32'd21076: dataIn1 = 32'd31
; 
32'd21077: dataIn1 = 32'd32
; 
32'd21078: dataIn1 = 32'd34
; 
32'd21079: dataIn1 = 32'd35
; 
32'd21080: dataIn1 = 32'd43
; 
32'd21081: dataIn1 = 32'd45
; 
32'd21082: dataIn1 = 32'd46
; 
32'd21083: dataIn1 = 32'd47
; 
32'd21084: dataIn1 = 32'd48
; 
32'd21085: dataIn1 = 32'd51
; 
32'd21086: dataIn1 = 32'd54
; 
32'd21087: dataIn1 = 32'd55
; 
32'd21088: dataIn1 = 32'd57
; 
32'd21089: dataIn1 = 32'd59
; 
32'd21090: dataIn1 = 32'd61
; 
32'd21091: dataIn1 = 32'd0
; 
32'd21092: dataIn1 = 32'd1
; 
32'd21093: dataIn1 = 32'd4
; 
32'd21094: dataIn1 = 32'd6
; 
32'd21095: dataIn1 = 32'd7
; 
32'd21096: dataIn1 = 32'd8
; 
32'd21097: dataIn1 = 32'd9
; 
32'd21098: dataIn1 = 32'd10
; 
32'd21099: dataIn1 = 32'd11
; 
32'd21100: dataIn1 = 32'd12
; 
32'd21101: dataIn1 = 32'd15
; 
32'd21102: dataIn1 = 32'd19
; 
32'd21103: dataIn1 = 32'd23
; 
32'd21104: dataIn1 = 32'd27
; 
32'd21105: dataIn1 = 32'd30
; 
32'd21106: dataIn1 = 32'd31
; 
32'd21107: dataIn1 = 32'd32
; 
32'd21108: dataIn1 = 32'd36
; 
32'd21109: dataIn1 = 32'd37
; 
32'd21110: dataIn1 = 32'd39
; 
32'd21111: dataIn1 = 32'd40
; 
32'd21112: dataIn1 = 32'd41
; 
32'd21113: dataIn1 = 32'd43
; 
32'd21114: dataIn1 = 32'd44
; 
32'd21115: dataIn1 = 32'd46
; 
32'd21116: dataIn1 = 32'd49
; 
32'd21117: dataIn1 = 32'd51
; 
32'd21118: dataIn1 = 32'd52
; 
32'd21119: dataIn1 = 32'd56
; 
32'd21120: dataIn1 = 32'd58
; 
32'd21121: dataIn1 = 32'd60
; 
32'd21122: dataIn1 = 32'd3
; 
32'd21123: dataIn1 = 32'd4
; 
32'd21124: dataIn1 = 32'd8
; 
32'd21125: dataIn1 = 32'd12
; 
32'd21126: dataIn1 = 32'd13
; 
32'd21127: dataIn1 = 32'd14
; 
32'd21128: dataIn1 = 32'd16
; 
32'd21129: dataIn1 = 32'd21
; 
32'd21130: dataIn1 = 32'd23
; 
32'd21131: dataIn1 = 32'd25
; 
32'd21132: dataIn1 = 32'd26
; 
32'd21133: dataIn1 = 32'd28
; 
32'd21134: dataIn1 = 32'd33
; 
32'd21135: dataIn1 = 32'd35
; 
32'd21136: dataIn1 = 32'd36
; 
32'd21137: dataIn1 = 32'd38
; 
32'd21138: dataIn1 = 32'd42
; 
32'd21139: dataIn1 = 32'd43
; 
32'd21140: dataIn1 = 32'd44
; 
32'd21141: dataIn1 = 32'd48
; 
32'd21142: dataIn1 = 32'd49
; 
32'd21143: dataIn1 = 32'd51
; 
32'd21144: dataIn1 = 32'd53
; 
32'd21145: dataIn1 = 32'd55
; 
32'd21146: dataIn1 = 32'd57
; 
32'd21147: dataIn1 = 32'd58
; 
32'd21148: dataIn1 = 32'd59
; 
32'd21149: dataIn1 = 32'd61
; 
32'd21150: dataIn1 = 32'd1
; 
32'd21151: dataIn1 = 32'd2
; 
32'd21152: dataIn1 = 32'd3
; 
32'd21153: dataIn1 = 32'd6
; 
32'd21154: dataIn1 = 32'd8
; 
32'd21155: dataIn1 = 32'd10
; 
32'd21156: dataIn1 = 32'd16
; 
32'd21157: dataIn1 = 32'd17
; 
32'd21158: dataIn1 = 32'd18
; 
32'd21159: dataIn1 = 32'd20
; 
32'd21160: dataIn1 = 32'd21
; 
32'd21161: dataIn1 = 32'd25
; 
32'd21162: dataIn1 = 32'd29
; 
32'd21163: dataIn1 = 32'd33
; 
32'd21164: dataIn1 = 32'd39
; 
32'd21165: dataIn1 = 32'd40
; 
32'd21166: dataIn1 = 32'd42
; 
32'd21167: dataIn1 = 32'd43
; 
32'd21168: dataIn1 = 32'd44
; 
32'd21169: dataIn1 = 32'd45
; 
32'd21170: dataIn1 = 32'd47
; 
32'd21171: dataIn1 = 32'd48
; 
32'd21172: dataIn1 = 32'd49
; 
32'd21173: dataIn1 = 32'd54
; 
32'd21174: dataIn1 = 32'd55
; 
32'd21175: dataIn1 = 32'd63
; 
32'd21176: dataIn1 = 32'd0
; 
32'd21177: dataIn1 = 32'd1
; 
32'd21178: dataIn1 = 32'd2
; 
32'd21179: dataIn1 = 32'd3
; 
32'd21180: dataIn1 = 32'd12
; 
32'd21181: dataIn1 = 32'd15
; 
32'd21182: dataIn1 = 32'd18
; 
32'd21183: dataIn1 = 32'd19
; 
32'd21184: dataIn1 = 32'd22
; 
32'd21185: dataIn1 = 32'd23
; 
32'd21186: dataIn1 = 32'd24
; 
32'd21187: dataIn1 = 32'd26
; 
32'd21188: dataIn1 = 32'd33
; 
32'd21189: dataIn1 = 32'd34
; 
32'd21190: dataIn1 = 32'd41
; 
32'd21191: dataIn1 = 32'd42
; 
32'd21192: dataIn1 = 32'd45
; 
32'd21193: dataIn1 = 32'd47
; 
32'd21194: dataIn1 = 32'd48
; 
32'd21195: dataIn1 = 32'd49
; 
32'd21196: dataIn1 = 32'd51
; 
32'd21197: dataIn1 = 32'd53
; 
32'd21198: dataIn1 = 32'd56
; 
32'd21199: dataIn1 = 32'd57
; 
32'd21200: dataIn1 = 32'd62
; 
32'd21201: dataIn1 = 32'd63
; 
32'd21202: dataIn1 = 32'd0
; 
32'd21203: dataIn1 = 32'd1
; 
32'd21204: dataIn1 = 32'd3
; 
32'd21205: dataIn1 = 32'd5
; 
32'd21206: dataIn1 = 32'd6
; 
32'd21207: dataIn1 = 32'd8
; 
32'd21208: dataIn1 = 32'd10
; 
32'd21209: dataIn1 = 32'd11
; 
32'd21210: dataIn1 = 32'd12
; 
32'd21211: dataIn1 = 32'd13
; 
32'd21212: dataIn1 = 32'd14
; 
32'd21213: dataIn1 = 32'd17
; 
32'd21214: dataIn1 = 32'd24
; 
32'd21215: dataIn1 = 32'd31
; 
32'd21216: dataIn1 = 32'd37
; 
32'd21217: dataIn1 = 32'd38
; 
32'd21218: dataIn1 = 32'd39
; 
32'd21219: dataIn1 = 32'd42
; 
32'd21220: dataIn1 = 32'd43
; 
32'd21221: dataIn1 = 32'd45
; 
32'd21222: dataIn1 = 32'd51
; 
32'd21223: dataIn1 = 32'd56
; 
32'd21224: dataIn1 = 32'd57
; 
32'd21225: dataIn1 = 32'd61
; 
32'd21226: dataIn1 = 32'd5
; 
32'd21227: dataIn1 = 32'd7
; 
32'd21228: dataIn1 = 32'd9
; 
32'd21229: dataIn1 = 32'd10
; 
32'd21230: dataIn1 = 32'd12
; 
32'd21231: dataIn1 = 32'd13
; 
32'd21232: dataIn1 = 32'd16
; 
32'd21233: dataIn1 = 32'd17
; 
32'd21234: dataIn1 = 32'd19
; 
32'd21235: dataIn1 = 32'd20
; 
32'd21236: dataIn1 = 32'd23
; 
32'd21237: dataIn1 = 32'd29
; 
32'd21238: dataIn1 = 32'd31
; 
32'd21239: dataIn1 = 32'd32
; 
32'd21240: dataIn1 = 32'd33
; 
32'd21241: dataIn1 = 32'd37
; 
32'd21242: dataIn1 = 32'd42
; 
32'd21243: dataIn1 = 32'd43
; 
32'd21244: dataIn1 = 32'd48
; 
32'd21245: dataIn1 = 32'd51
; 
32'd21246: dataIn1 = 32'd52
; 
32'd21247: dataIn1 = 32'd54
; 
32'd21248: dataIn1 = 32'd4
; 
32'd21249: dataIn1 = 32'd6
; 
32'd21250: dataIn1 = 32'd9
; 
32'd21251: dataIn1 = 32'd13
; 
32'd21252: dataIn1 = 32'd16
; 
32'd21253: dataIn1 = 32'd19
; 
32'd21254: dataIn1 = 32'd23
; 
32'd21255: dataIn1 = 32'd29
; 
32'd21256: dataIn1 = 32'd32
; 
32'd21257: dataIn1 = 32'd34
; 
32'd21258: dataIn1 = 32'd39
; 
32'd21259: dataIn1 = 32'd40
; 
32'd21260: dataIn1 = 32'd49
; 
32'd21261: dataIn1 = 32'd51
; 
32'd21262: dataIn1 = 32'd52
; 
32'd21263: dataIn1 = 32'd55
; 
32'd21264: dataIn1 = 32'd57
; 
32'd21265: dataIn1 = 32'd59
; 
32'd21266: dataIn1 = 32'd60
; 
32'd21267: dataIn1 = 32'd13
; 
32'd21268: dataIn1 = 32'd17
; 
32'd21269: dataIn1 = 32'd20
; 
32'd21270: dataIn1 = 32'd22
; 
32'd21271: dataIn1 = 32'd25
; 
32'd21272: dataIn1 = 32'd26
; 
32'd21273: dataIn1 = 32'd30
; 
32'd21274: dataIn1 = 32'd33
; 
32'd21275: dataIn1 = 32'd35
; 
32'd21276: dataIn1 = 32'd36
; 
32'd21277: dataIn1 = 32'd44
; 
32'd21278: dataIn1 = 32'd45
; 
32'd21279: dataIn1 = 32'd46
; 
32'd21280: dataIn1 = 32'd48
; 
32'd21281: dataIn1 = 32'd49
; 
32'd21282: dataIn1 = 32'd51
; 
32'd21283: dataIn1 = 32'd53
; 
32'd21284: dataIn1 = 32'd54
; 
32'd21285: dataIn1 = 32'd55
; 
32'd21286: dataIn1 = 32'd62
; 
32'd21287: dataIn1 = 32'd63
; 
32'd21288: dataIn1 = 32'd5
; 
32'd21289: dataIn1 = 32'd6
; 
32'd21290: dataIn1 = 32'd11
; 
32'd21291: dataIn1 = 32'd12
; 
32'd21292: dataIn1 = 32'd25
; 
32'd21293: dataIn1 = 32'd28
; 
32'd21294: dataIn1 = 32'd40
; 
32'd21295: dataIn1 = 32'd41
; 
32'd21296: dataIn1 = 32'd44
; 
32'd21297: dataIn1 = 32'd47
; 
32'd21298: dataIn1 = 32'd57
; 
32'd21299: dataIn1 = 32'd58
; 
32'd21300: dataIn1 = 32'd59
; 
32'd21301: dataIn1 = 32'd62
; 
32'd21302: dataIn1 = 32'd; 
32'd21303: dataIn1 = 32'd; 
32'd21304: dataIn1 = 32'd; 
32'd21305: dataIn1 = 32'd; 
32'd21306: dataIn1 = 32'd; 
32'd21307: dataIn1 = 32'd; 
32'd21308: dataIn1 = 32'd; 
32'd21309: dataIn1 = 32'd; 
32'd21310: dataIn1 = 32'd; 
32'd21311: dataIn1 = 32'd; 
32'd21312: dataIn1 = 32'd; 
32'd21313: dataIn1 = 32'd; 
32'd21314: dataIn1 = 32'd; 
32'd21315: dataIn1 = 32'd; 
32'd21316: dataIn1 = 32'd; 
32'd21317: dataIn1 = 32'd; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd14; 
32'd3: dataIn2 = 32'd73; 
32'd4: dataIn2 = 32'd42; 
32'd5: dataIn2 = 32'd100; 
32'd6: dataIn2 = 32'd15; 
32'd7: dataIn2 = 32'd53; 
32'd8: dataIn2 = 32'd68; 
32'd9: dataIn2 = 32'd56; 
32'd10: dataIn2 = 32'd57; 
32'd11: dataIn2 = 32'd92; 
32'd12: dataIn2 = 32'd10; 
32'd13: dataIn2 = 32'd52; 
32'd14: dataIn2 = 32'd99; 
32'd15: dataIn2 = 32'd99; 
32'd16: dataIn2 = 32'd64; 
32'd17: dataIn2 = 32'd6; 
32'd18: dataIn2 = 32'd77; 
32'd19: dataIn2 = 32'd80; 
32'd20: dataIn2 = 32'd29; 
32'd21: dataIn2 = 32'd71; 
32'd22: dataIn2 = 32'd100; 
32'd23: dataIn2 = 32'd34; 
32'd24: dataIn2 = 32'd32; 
32'd25: dataIn2 = 32'd25; 
32'd26: dataIn2 = 32'd23; 
32'd27: dataIn2 = 32'd46; 
32'd28: dataIn2 = 32'd72; 
32'd29: dataIn2 = 32'd76; 
32'd30: dataIn2 = 32'd85; 
32'd31: dataIn2 = 32'd59; 
32'd32: dataIn2 = 32'd42; 
32'd33: dataIn2 = 32'd36; 
32'd34: dataIn2 = 32'd65; 
32'd35: dataIn2 = 32'd42; 
32'd36: dataIn2 = 32'd23; 
32'd37: dataIn2 = 32'd84; 
32'd38: dataIn2 = 32'd40; 
32'd39: dataIn2 = 32'd59; 
32'd40: dataIn2 = 32'd85; 
32'd41: dataIn2 = 32'd28; 
32'd42: dataIn2 = 32'd35; 
32'd43: dataIn2 = 32'd14; 
32'd44: dataIn2 = 32'd37; 
32'd45: dataIn2 = 32'd97; 
32'd46: dataIn2 = 32'd3; 
32'd47: dataIn2 = 32'd70; 
32'd48: dataIn2 = 32'd74; 
32'd49: dataIn2 = 32'd2; 
32'd50: dataIn2 = 32'd24; 
32'd51: dataIn2 = 32'd22; 
32'd52: dataIn2 = 32'd39; 
32'd53: dataIn2 = 32'd89; 
32'd54: dataIn2 = 32'd46; 
32'd55: dataIn2 = 32'd99; 
32'd56: dataIn2 = 32'd45; 
32'd57: dataIn2 = 32'd27; 
32'd58: dataIn2 = 32'd85; 
32'd59: dataIn2 = 32'd56; 
32'd60: dataIn2 = 32'd90; 
32'd61: dataIn2 = 32'd61; 
32'd62: dataIn2 = 32'd80; 
32'd63: dataIn2 = 32'd7; 
32'd64: dataIn2 = 32'd28; 
32'd65: dataIn2 = 32'd69; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd330: dataIn2 = 32'd10; 
32'd331: dataIn2 = 32'd20; 
32'd332: dataIn2 = 32'd34; 
32'd333: dataIn2 = 32'd99; 
32'd334: dataIn2 = 32'd59; 
32'd335: dataIn2 = 32'd1; 
32'd336: dataIn2 = 32'd8; 
32'd337: dataIn2 = 32'd55; 
32'd338: dataIn2 = 32'd34; 
32'd339: dataIn2 = 32'd3; 
32'd340: dataIn2 = 32'd92; 
32'd341: dataIn2 = 32'd83; 
32'd342: dataIn2 = 32'd80; 
32'd343: dataIn2 = 32'd77; 
32'd344: dataIn2 = 32'd38; 
32'd345: dataIn2 = 32'd80; 
32'd346: dataIn2 = 32'd88; 
32'd347: dataIn2 = 32'd20; 
32'd348: dataIn2 = 32'd19; 
32'd349: dataIn2 = 32'd12; 
32'd350: dataIn2 = 32'd73; 
32'd351: dataIn2 = 32'd98; 
32'd352: dataIn2 = 32'd65; 
32'd353: dataIn2 = 32'd44; 
32'd354: dataIn2 = 32'd74; 
32'd355: dataIn2 = 32'd73; 
32'd356: dataIn2 = 32'd43; 
32'd357: dataIn2 = 32'd91; 
32'd358: dataIn2 = 32'd45; 
32'd359: dataIn2 = 32'd54; 
32'd360: dataIn2 = 32'd61; 
32'd361: dataIn2 = 32'd87; 
32'd362: dataIn2 = 32'd2; 
32'd363: dataIn2 = 32'd59; 
32'd364: dataIn2 = 32'd62; 
32'd365: dataIn2 = 32'd21; 
32'd366: dataIn2 = 32'd96; 
32'd367: dataIn2 = 32'd44; 
32'd368: dataIn2 = 32'd23; 
32'd369: dataIn2 = 32'd91; 
32'd370: dataIn2 = 32'd16; 
32'd371: dataIn2 = 32'd65; 
32'd372: dataIn2 = 32'd98; 
32'd373: dataIn2 = 32'd92; 
32'd374: dataIn2 = 32'd85; 
32'd375: dataIn2 = 32'd89; 
32'd376: dataIn2 = 32'd67; 
32'd377: dataIn2 = 32'd79; 
32'd378: dataIn2 = 32'd67; 
32'd379: dataIn2 = 32'd99; 
32'd380: dataIn2 = 32'd82; 
32'd381: dataIn2 = 32'd32; 
32'd382: dataIn2 = 32'd13; 
32'd383: dataIn2 = 32'd91; 
32'd384: dataIn2 = 32'd47; 
32'd385: dataIn2 = 32'd91; 
32'd386: dataIn2 = 32'd9; 
32'd387: dataIn2 = 32'd32; 
32'd388: dataIn2 = 32'd48; 
32'd389: dataIn2 = 32'd11; 
32'd390: dataIn2 = 32'd8; 
32'd391: dataIn2 = 32'd30; 
32'd392: dataIn2 = 32'd98; 
32'd393: dataIn2 = 32'd98; 
32'd394: dataIn2 = 32'd12; 
32'd395: dataIn2 = 32'd27; 
32'd396: dataIn2 = 32'd46; 
32'd397: dataIn2 = 32'd18; 
32'd398: dataIn2 = 32'd71; 
32'd399: dataIn2 = 32'd62; 
32'd400: dataIn2 = 32'd57; 
32'd401: dataIn2 = 32'd34; 
32'd402: dataIn2 = 32'd43; 
32'd403: dataIn2 = 32'd0; 
32'd404: dataIn2 = 32'd49; 
32'd405: dataIn2 = 32'd64; 
32'd406: dataIn2 = 32'd69; 
32'd407: dataIn2 = 32'd55; 
32'd408: dataIn2 = 32'd38; 
32'd409: dataIn2 = 32'd18; 
32'd410: dataIn2 = 32'd12; 
32'd411: dataIn2 = 32'd21; 
32'd412: dataIn2 = 32'd1; 
32'd413: dataIn2 = 32'd79; 
32'd414: dataIn2 = 32'd99; 
32'd415: dataIn2 = 32'd78; 
32'd416: dataIn2 = 32'd80; 
32'd417: dataIn2 = 32'd51; 
32'd418: dataIn2 = 32'd48; 
32'd419: dataIn2 = 32'd55; 
32'd420: dataIn2 = 32'd81; 
32'd421: dataIn2 = 32'd62; 
32'd422: dataIn2 = 32'd31; 
32'd423: dataIn2 = 32'd25; 
32'd424: dataIn2 = 32'd76; 
32'd425: dataIn2 = 32'd21; 
32'd426: dataIn2 = 32'd9; 
32'd427: dataIn2 = 32'd85; 
32'd428: dataIn2 = 32'd81; 
32'd429: dataIn2 = 32'd32; 
32'd430: dataIn2 = 32'd4; 
32'd431: dataIn2 = 32'd4; 
32'd432: dataIn2 = 32'd14; 
32'd433: dataIn2 = 32'd94; 
32'd434: dataIn2 = 32'd12; 
32'd435: dataIn2 = 32'd35; 
32'd436: dataIn2 = 32'd93; 
32'd437: dataIn2 = 32'd76; 
32'd438: dataIn2 = 32'd95; 
32'd439: dataIn2 = 32'd8; 
32'd440: dataIn2 = 32'd9; 
32'd441: dataIn2 = 32'd91; 
32'd442: dataIn2 = 32'd69; 
32'd443: dataIn2 = 32'd5; 
32'd444: dataIn2 = 32'd32; 
32'd445: dataIn2 = 32'd46; 
32'd446: dataIn2 = 32'd96; 
32'd447: dataIn2 = 32'd28; 
32'd448: dataIn2 = 32'd20; 
32'd449: dataIn2 = 32'd59; 
32'd450: dataIn2 = 32'd89; 
32'd451: dataIn2 = 32'd11; 
32'd452: dataIn2 = 32'd55; 
32'd453: dataIn2 = 32'd57; 
32'd454: dataIn2 = 32'd93; 
32'd455: dataIn2 = 32'd63; 
32'd456: dataIn2 = 32'd56; 
32'd457: dataIn2 = 32'd42; 
32'd458: dataIn2 = 32'd3; 
32'd459: dataIn2 = 32'd93; 
32'd460: dataIn2 = 32'd60; 
32'd461: dataIn2 = 32'd5; 
32'd462: dataIn2 = 32'd28; 
32'd463: dataIn2 = 32'd65; 
32'd464: dataIn2 = 32'd41; 
32'd465: dataIn2 = 32'd71; 
32'd466: dataIn2 = 32'd54; 
32'd467: dataIn2 = 32'd94; 
32'd468: dataIn2 = 32'd25; 
32'd469: dataIn2 = 32'd57; 
32'd470: dataIn2 = 32'd17; 
32'd471: dataIn2 = 32'd82; 
32'd472: dataIn2 = 32'd99; 
32'd473: dataIn2 = 32'd98; 
32'd474: dataIn2 = 32'd14; 
32'd475: dataIn2 = 32'd3; 
32'd476: dataIn2 = 32'd8; 
32'd477: dataIn2 = 32'd82; 
32'd478: dataIn2 = 32'd99; 
32'd479: dataIn2 = 32'd18; 
32'd480: dataIn2 = 32'd83; 
32'd481: dataIn2 = 32'd59; 
32'd482: dataIn2 = 32'd46; 
32'd483: dataIn2 = 32'd38; 
32'd484: dataIn2 = 32'd38; 
32'd485: dataIn2 = 32'd56; 
32'd486: dataIn2 = 32'd55; 
32'd487: dataIn2 = 32'd5; 
32'd488: dataIn2 = 32'd64; 
32'd489: dataIn2 = 32'd71; 
32'd490: dataIn2 = 32'd73; 
32'd491: dataIn2 = 32'd6; 
32'd492: dataIn2 = 32'd91; 
32'd493: dataIn2 = 32'd46; 
32'd494: dataIn2 = 32'd30; 
32'd495: dataIn2 = 32'd57; 
32'd496: dataIn2 = 32'd26; 
32'd497: dataIn2 = 32'd29; 
32'd498: dataIn2 = 32'd89; 
32'd499: dataIn2 = 32'd23; 
32'd500: dataIn2 = 32'd66; 
32'd501: dataIn2 = 32'd50; 
32'd502: dataIn2 = 32'd14; 
32'd503: dataIn2 = 32'd58; 
32'd504: dataIn2 = 32'd24; 
32'd505: dataIn2 = 32'd34; 
32'd506: dataIn2 = 32'd50; 
32'd507: dataIn2 = 32'd36; 
32'd508: dataIn2 = 32'd63; 
32'd509: dataIn2 = 32'd30; 
32'd510: dataIn2 = 32'd25; 
32'd511: dataIn2 = 32'd43; 
32'd512: dataIn2 = 32'd22; 
32'd513: dataIn2 = 32'd39; 
32'd514: dataIn2 = 32'd20; 
32'd515: dataIn2 = 32'd91; 
32'd516: dataIn2 = 32'd83; 
32'd517: dataIn2 = 32'd90; 
32'd518: dataIn2 = 32'd84; 
32'd519: dataIn2 = 32'd53; 
32'd520: dataIn2 = 32'd41; 
32'd521: dataIn2 = 32'd39; 
32'd522: dataIn2 = 32'd63; 
32'd523: dataIn2 = 32'd90; 
32'd524: dataIn2 = 32'd70; 
32'd525: dataIn2 = 32'd83; 
32'd526: dataIn2 = 32'd12; 
32'd527: dataIn2 = 32'd47; 
32'd528: dataIn2 = 32'd9; 
32'd529: dataIn2 = 32'd50; 
32'd530: dataIn2 = 32'd94; 
32'd531: dataIn2 = 32'd58; 
32'd532: dataIn2 = 32'd14; 
32'd533: dataIn2 = 32'd42; 
32'd534: dataIn2 = 32'd6; 
32'd535: dataIn2 = 32'd7; 
32'd536: dataIn2 = 32'd5; 
32'd537: dataIn2 = 32'd31; 
32'd538: dataIn2 = 32'd65; 
32'd539: dataIn2 = 32'd96; 
32'd540: dataIn2 = 32'd93; 
32'd541: dataIn2 = 32'd26; 
32'd542: dataIn2 = 32'd46; 
32'd543: dataIn2 = 32'd32; 
32'd544: dataIn2 = 32'd48; 
32'd545: dataIn2 = 32'd63; 
32'd546: dataIn2 = 32'd22; 
32'd547: dataIn2 = 32'd18; 
32'd548: dataIn2 = 32'd53; 
32'd549: dataIn2 = 32'd79; 
32'd550: dataIn2 = 32'd18; 
32'd551: dataIn2 = 32'd67; 
32'd552: dataIn2 = 32'd25; 
32'd553: dataIn2 = 32'd16; 
32'd554: dataIn2 = 32'd40; 
32'd555: dataIn2 = 32'd56; 
32'd556: dataIn2 = 32'd80; 
32'd557: dataIn2 = 32'd31; 
32'd558: dataIn2 = 32'd58; 
32'd559: dataIn2 = 32'd25; 
32'd560: dataIn2 = 32'd94; 
32'd561: dataIn2 = 32'd43; 
32'd562: dataIn2 = 32'd43; 
32'd563: dataIn2 = 32'd91; 
32'd564: dataIn2 = 32'd36; 
32'd565: dataIn2 = 32'd63; 
32'd566: dataIn2 = 32'd55; 
32'd567: dataIn2 = 32'd97; 
32'd568: dataIn2 = 32'd75; 
32'd569: dataIn2 = 32'd83; 
32'd570: dataIn2 = 32'd81; 
32'd571: dataIn2 = 32'd52; 
32'd572: dataIn2 = 32'd10; 
32'd573: dataIn2 = 32'd5; 
32'd574: dataIn2 = 32'd13; 
32'd575: dataIn2 = 32'd53; 
32'd576: dataIn2 = 32'd64; 
32'd577: dataIn2 = 32'd70; 
32'd578: dataIn2 = 32'd26; 
32'd579: dataIn2 = 32'd85; 
32'd580: dataIn2 = 32'd34; 
32'd581: dataIn2 = 32'd94; 
32'd582: dataIn2 = 32'd15; 
32'd583: dataIn2 = 32'd20; 
32'd584: dataIn2 = 32'd43; 
32'd585: dataIn2 = 32'd65; 
32'd586: dataIn2 = 32'd98; 
32'd587: dataIn2 = 32'd51; 
32'd588: dataIn2 = 32'd65; 
32'd589: dataIn2 = 32'd24; 
32'd590: dataIn2 = 32'd34; 
32'd591: dataIn2 = 32'd38; 
32'd592: dataIn2 = 32'd59; 
32'd593: dataIn2 = 32'd37; 
32'd594: dataIn2 = 32'd15; 
32'd595: dataIn2 = 32'd25; 
32'd596: dataIn2 = 32'd4; 
32'd597: dataIn2 = 32'd17; 
32'd598: dataIn2 = 32'd52; 
32'd599: dataIn2 = 32'd0; 
32'd600: dataIn2 = 32'd26; 
32'd601: dataIn2 = 32'd68; 
32'd602: dataIn2 = 32'd20; 
32'd603: dataIn2 = 32'd32; 
32'd604: dataIn2 = 32'd92; 
32'd605: dataIn2 = 32'd24; 
32'd606: dataIn2 = 32'd92; 
32'd607: dataIn2 = 32'd18; 
32'd608: dataIn2 = 32'd82; 
32'd609: dataIn2 = 32'd51; 
32'd610: dataIn2 = 32'd65; 
32'd611: dataIn2 = 32'd4; 
32'd612: dataIn2 = 32'd46; 
32'd613: dataIn2 = 32'd0; 
32'd614: dataIn2 = 32'd86; 
32'd615: dataIn2 = 32'd51; 
32'd616: dataIn2 = 32'd60; 
32'd617: dataIn2 = 32'd76; 
32'd618: dataIn2 = 32'd78; 
32'd619: dataIn2 = 32'd86; 
32'd620: dataIn2 = 32'd68; 
32'd621: dataIn2 = 32'd60; 
32'd622: dataIn2 = 32'd77; 
32'd623: dataIn2 = 32'd3; 
32'd624: dataIn2 = 32'd11; 
32'd625: dataIn2 = 32'd71; 
32'd626: dataIn2 = 32'd63; 
32'd627: dataIn2 = 32'd55; 
32'd628: dataIn2 = 32'd7; 
32'd629: dataIn2 = 32'd2; 
32'd630: dataIn2 = 32'd12; 
32'd631: dataIn2 = 32'd91; 
32'd632: dataIn2 = 32'd92; 
32'd633: dataIn2 = 32'd44; 
32'd634: dataIn2 = 32'd60; 
32'd635: dataIn2 = 32'd91; 
32'd636: dataIn2 = 32'd57; 
32'd637: dataIn2 = 32'd24; 
32'd638: dataIn2 = 32'd56; 
32'd639: dataIn2 = 32'd10; 
32'd640: dataIn2 = 32'd20; 
32'd641: dataIn2 = 32'd13; 
32'd642: dataIn2 = 32'd64; 
32'd643: dataIn2 = 32'd5; 
32'd644: dataIn2 = 32'd28; 
32'd645: dataIn2 = 32'd51; 
32'd646: dataIn2 = 32'd89; 
32'd647: dataIn2 = 32'd8; 
32'd648: dataIn2 = 32'd87; 
32'd649: dataIn2 = 32'd68; 
32'd650: dataIn2 = 32'd21; 
32'd651: dataIn2 = 32'd39; 
32'd652: dataIn2 = 32'd60; 
32'd653: dataIn2 = 32'd10; 
32'd654: dataIn2 = 32'd39; 
32'd655: dataIn2 = 32'd55; 
32'd656: dataIn2 = 32'd67; 
32'd657: dataIn2 = 32'd88; 
32'd658: dataIn2 = 32'd1; 
32'd659: dataIn2 = 32'd18; 
32'd660: dataIn2 = 32'd64; 
32'd661: dataIn2 = 32'd93; 
32'd662: dataIn2 = 32'd43; 
32'd663: dataIn2 = 32'd30; 
32'd664: dataIn2 = 32'd7; 
32'd665: dataIn2 = 32'd29; 
32'd666: dataIn2 = 32'd68; 
32'd667: dataIn2 = 32'd26; 
32'd668: dataIn2 = 32'd54; 
32'd669: dataIn2 = 32'd48; 
32'd670: dataIn2 = 32'd14; 
32'd671: dataIn2 = 32'd78; 
32'd672: dataIn2 = 32'd84; 
32'd673: dataIn2 = 32'd73; 
32'd674: dataIn2 = 32'd71; 
32'd675: dataIn2 = 32'd33; 
32'd676: dataIn2 = 32'd31; 
32'd677: dataIn2 = 32'd38; 
32'd678: dataIn2 = 32'd52; 
32'd679: dataIn2 = 32'd62; 
32'd680: dataIn2 = 32'd0; 
32'd681: dataIn2 = 32'd87; 
32'd682: dataIn2 = 32'd43; 
32'd683: dataIn2 = 32'd82; 
32'd684: dataIn2 = 32'd3; 
32'd685: dataIn2 = 32'd83; 
32'd686: dataIn2 = 32'd34; 
32'd687: dataIn2 = 32'd13; 
32'd688: dataIn2 = 32'd1; 
32'd689: dataIn2 = 32'd30; 
32'd690: dataIn2 = 32'd89; 
32'd691: dataIn2 = 32'd97; 
32'd692: dataIn2 = 32'd78; 
32'd693: dataIn2 = 32'd66; 
32'd694: dataIn2 = 32'd27; 
32'd695: dataIn2 = 32'd53; 
32'd696: dataIn2 = 32'd70; 
32'd697: dataIn2 = 32'd99; 
32'd698: dataIn2 = 32'd29; 
32'd699: dataIn2 = 32'd90; 
32'd700: dataIn2 = 32'd39; 
32'd701: dataIn2 = 32'd99; 
32'd702: dataIn2 = 32'd55; 
32'd703: dataIn2 = 32'd38; 
32'd704: dataIn2 = 32'd70; 
32'd705: dataIn2 = 32'd25; 
32'd706: dataIn2 = 32'd69; 
32'd707: dataIn2 = 32'd70; 
32'd708: dataIn2 = 32'd29; 
32'd709: dataIn2 = 32'd95; 
32'd710: dataIn2 = 32'd38; 
32'd711: dataIn2 = 32'd51; 
32'd712: dataIn2 = 32'd86; 
32'd713: dataIn2 = 32'd1; 
32'd714: dataIn2 = 32'd24; 
32'd715: dataIn2 = 32'd77; 
32'd716: dataIn2 = 32'd98; 
32'd717: dataIn2 = 32'd35; 
32'd718: dataIn2 = 32'd12; 
32'd719: dataIn2 = 32'd14; 
32'd720: dataIn2 = 32'd82; 
32'd721: dataIn2 = 32'd72; 
32'd722: dataIn2 = 32'd82; 
32'd723: dataIn2 = 32'd72; 
32'd724: dataIn2 = 32'd87; 
32'd725: dataIn2 = 32'd25; 
32'd726: dataIn2 = 32'd24; 
32'd727: dataIn2 = 32'd2; 
32'd728: dataIn2 = 32'd71; 
32'd729: dataIn2 = 32'd93; 
32'd730: dataIn2 = 32'd55; 
32'd731: dataIn2 = 32'd95; 
32'd732: dataIn2 = 32'd42; 
32'd733: dataIn2 = 32'd87; 
32'd734: dataIn2 = 32'd0; 
32'd735: dataIn2 = 32'd8; 
32'd736: dataIn2 = 32'd12; 
32'd737: dataIn2 = 32'd67; 
32'd738: dataIn2 = 32'd31; 
32'd739: dataIn2 = 32'd53; 
32'd740: dataIn2 = 32'd30; 
32'd741: dataIn2 = 32'd44; 
32'd742: dataIn2 = 32'd47; 
32'd743: dataIn2 = 32'd28; 
32'd744: dataIn2 = 32'd83; 
32'd745: dataIn2 = 32'd100; 
32'd746: dataIn2 = 32'd1; 
32'd747: dataIn2 = 32'd23; 
32'd748: dataIn2 = 32'd18; 
32'd749: dataIn2 = 32'd45; 
32'd750: dataIn2 = 32'd69; 
32'd751: dataIn2 = 32'd98; 
32'd752: dataIn2 = 32'd99; 
32'd753: dataIn2 = 32'd75; 
32'd754: dataIn2 = 32'd70; 
32'd755: dataIn2 = 32'd35; 
32'd756: dataIn2 = 32'd44; 
32'd757: dataIn2 = 32'd96; 
32'd758: dataIn2 = 32'd30; 
32'd759: dataIn2 = 32'd44; 
32'd760: dataIn2 = 32'd14; 
32'd761: dataIn2 = 32'd53; 
32'd762: dataIn2 = 32'd89; 
32'd763: dataIn2 = 32'd42; 
32'd764: dataIn2 = 32'd12; 
32'd765: dataIn2 = 32'd18; 
32'd766: dataIn2 = 32'd23; 
32'd767: dataIn2 = 32'd36; 
32'd768: dataIn2 = 32'd2; 
32'd769: dataIn2 = 32'd62; 
32'd770: dataIn2 = 32'd86; 
32'd771: dataIn2 = 32'd29; 
32'd772: dataIn2 = 32'd20; 
32'd773: dataIn2 = 32'd74; 
32'd774: dataIn2 = 32'd11; 
32'd775: dataIn2 = 32'd44; 
32'd776: dataIn2 = 32'd55; 
32'd777: dataIn2 = 32'd53; 
32'd778: dataIn2 = 32'd82; 
32'd779: dataIn2 = 32'd50; 
32'd780: dataIn2 = 32'd2; 
32'd781: dataIn2 = 32'd66; 
32'd782: dataIn2 = 32'd98; 
32'd783: dataIn2 = 32'd39; 
32'd784: dataIn2 = 32'd89; 
32'd785: dataIn2 = 32'd85; 
32'd786: dataIn2 = 32'd41; 
32'd787: dataIn2 = 32'd95; 
32'd788: dataIn2 = 32'd78; 
32'd789: dataIn2 = 32'd62; 
32'd790: dataIn2 = 32'd23; 
32'd791: dataIn2 = 32'd64; 
32'd792: dataIn2 = 32'd20; 
32'd793: dataIn2 = 32'd88; 
32'd794: dataIn2 = 32'd47; 
32'd795: dataIn2 = 32'd25; 
32'd796: dataIn2 = 32'd70; 
32'd797: dataIn2 = 32'd90; 
32'd798: dataIn2 = 32'd86; 
32'd799: dataIn2 = 32'd56; 
32'd800: dataIn2 = 32'd17; 
32'd801: dataIn2 = 32'd74; 
32'd802: dataIn2 = 32'd10; 
32'd803: dataIn2 = 32'd31; 
32'd804: dataIn2 = 32'd27; 
32'd805: dataIn2 = 32'd42; 
32'd806: dataIn2 = 32'd91; 
32'd807: dataIn2 = 32'd25; 
32'd808: dataIn2 = 32'd17; 
32'd809: dataIn2 = 32'd57; 
32'd810: dataIn2 = 32'd69; 
32'd811: dataIn2 = 32'd83; 
32'd812: dataIn2 = 32'd85; 
32'd813: dataIn2 = 32'd72; 
32'd814: dataIn2 = 32'd18; 
32'd815: dataIn2 = 32'd24; 
32'd816: dataIn2 = 32'd11; 
32'd817: dataIn2 = 32'd17; 
32'd818: dataIn2 = 32'd10; 
32'd819: dataIn2 = 32'd39; 
32'd820: dataIn2 = 32'd59; 
32'd821: dataIn2 = 32'd27; 
32'd822: dataIn2 = 32'd65; 
32'd823: dataIn2 = 32'd61; 
32'd824: dataIn2 = 32'd9; 
32'd825: dataIn2 = 32'd47; 
32'd826: dataIn2 = 32'd89; 
32'd827: dataIn2 = 32'd7; 
32'd828: dataIn2 = 32'd0; 
32'd829: dataIn2 = 32'd31; 
32'd830: dataIn2 = 32'd20; 
32'd831: dataIn2 = 32'd99; 
32'd832: dataIn2 = 32'd90; 
32'd833: dataIn2 = 32'd86; 
32'd834: dataIn2 = 32'd99; 
32'd835: dataIn2 = 32'd90; 
32'd836: dataIn2 = 32'd2; 
32'd837: dataIn2 = 32'd79; 
32'd838: dataIn2 = 32'd48; 
32'd839: dataIn2 = 32'd0; 
32'd840: dataIn2 = 32'd20; 
32'd841: dataIn2 = 32'd8; 
32'd842: dataIn2 = 32'd34; 
32'd843: dataIn2 = 32'd21; 
32'd844: dataIn2 = 32'd69; 
32'd845: dataIn2 = 32'd10; 
32'd846: dataIn2 = 32'd38; 
32'd847: dataIn2 = 32'd99; 
32'd848: dataIn2 = 32'd19; 
32'd849: dataIn2 = 32'd54; 
32'd850: dataIn2 = 32'd47; 
32'd851: dataIn2 = 32'd59; 
32'd852: dataIn2 = 32'd22; 
32'd853: dataIn2 = 32'd24; 
32'd854: dataIn2 = 32'd37; 
32'd855: dataIn2 = 32'd74; 
32'd856: dataIn2 = 32'd77; 
32'd857: dataIn2 = 32'd8; 
32'd858: dataIn2 = 32'd1; 
32'd859: dataIn2 = 32'd13; 
32'd860: dataIn2 = 32'd12; 
32'd861: dataIn2 = 32'd19; 
32'd862: dataIn2 = 32'd96; 
32'd863: dataIn2 = 32'd48; 
32'd864: dataIn2 = 32'd40; 
32'd865: dataIn2 = 32'd9; 
32'd866: dataIn2 = 32'd97; 
32'd867: dataIn2 = 32'd24; 
32'd868: dataIn2 = 32'd9; 
32'd869: dataIn2 = 32'd98; 
32'd870: dataIn2 = 32'd99; 
32'd871: dataIn2 = 32'd14; 
32'd872: dataIn2 = 32'd60; 
32'd873: dataIn2 = 32'd25; 
32'd874: dataIn2 = 32'd11; 
32'd875: dataIn2 = 32'd96; 
32'd876: dataIn2 = 32'd63; 
32'd877: dataIn2 = 32'd75; 
32'd878: dataIn2 = 32'd97; 
32'd879: dataIn2 = 32'd39; 
32'd880: dataIn2 = 32'd93; 
32'd881: dataIn2 = 32'd97; 
32'd882: dataIn2 = 32'd14; 
32'd883: dataIn2 = 32'd11; 
32'd884: dataIn2 = 32'd7; 
32'd885: dataIn2 = 32'd57; 
32'd886: dataIn2 = 32'd100; 
32'd887: dataIn2 = 32'd50; 
32'd888: dataIn2 = 32'd14; 
32'd889: dataIn2 = 32'd72; 
32'd890: dataIn2 = 32'd22; 
32'd891: dataIn2 = 32'd71; 
32'd892: dataIn2 = 32'd83; 
32'd893: dataIn2 = 32'd43; 
32'd894: dataIn2 = 32'd10; 
32'd895: dataIn2 = 32'd87; 
32'd896: dataIn2 = 32'd42; 
32'd897: dataIn2 = 32'd31; 
32'd898: dataIn2 = 32'd8; 
32'd899: dataIn2 = 32'd81; 
32'd900: dataIn2 = 32'd28; 
32'd901: dataIn2 = 32'd69; 
32'd902: dataIn2 = 32'd37; 
32'd903: dataIn2 = 32'd55; 
32'd904: dataIn2 = 32'd5; 
32'd905: dataIn2 = 32'd99; 
32'd906: dataIn2 = 32'd81; 
32'd907: dataIn2 = 32'd32; 
32'd908: dataIn2 = 32'd16; 
32'd909: dataIn2 = 32'd84; 
32'd910: dataIn2 = 32'd13; 
32'd911: dataIn2 = 32'd6; 
32'd912: dataIn2 = 32'd60; 
32'd913: dataIn2 = 32'd8; 
32'd914: dataIn2 = 32'd92; 
32'd915: dataIn2 = 32'd12; 
32'd916: dataIn2 = 32'd98; 
32'd917: dataIn2 = 32'd58; 
32'd918: dataIn2 = 32'd73; 
32'd919: dataIn2 = 32'd17; 
32'd920: dataIn2 = 32'd29; 
32'd921: dataIn2 = 32'd83; 
32'd922: dataIn2 = 32'd53; 
32'd923: dataIn2 = 32'd36; 
32'd924: dataIn2 = 32'd82; 
32'd925: dataIn2 = 32'd57; 
32'd926: dataIn2 = 32'd70; 
32'd927: dataIn2 = 32'd10; 
32'd928: dataIn2 = 32'd53; 
32'd929: dataIn2 = 32'd96; 
32'd930: dataIn2 = 32'd80; 
32'd931: dataIn2 = 32'd34; 
32'd932: dataIn2 = 32'd82; 
32'd933: dataIn2 = 32'd40; 
32'd934: dataIn2 = 32'd67; 
32'd935: dataIn2 = 32'd54; 
32'd936: dataIn2 = 32'd29; 
32'd937: dataIn2 = 32'd72; 
32'd938: dataIn2 = 32'd95; 
32'd939: dataIn2 = 32'd28; 
32'd940: dataIn2 = 32'd45; 
32'd941: dataIn2 = 32'd99; 
32'd942: dataIn2 = 32'd14; 
32'd943: dataIn2 = 32'd68; 
32'd944: dataIn2 = 32'd94; 
32'd945: dataIn2 = 32'd51; 
32'd946: dataIn2 = 32'd20; 
32'd947: dataIn2 = 32'd1; 
32'd948: dataIn2 = 32'd41; 
32'd949: dataIn2 = 32'd65; 
32'd950: dataIn2 = 32'd78; 
32'd951: dataIn2 = 32'd34; 
32'd952: dataIn2 = 32'd8; 
32'd953: dataIn2 = 32'd23; 
32'd954: dataIn2 = 32'd92; 
32'd955: dataIn2 = 32'd62; 
32'd956: dataIn2 = 32'd73; 
32'd957: dataIn2 = 32'd22; 
32'd958: dataIn2 = 32'd62; 
32'd959: dataIn2 = 32'd35; 
32'd960: dataIn2 = 32'd56; 
32'd961: dataIn2 = 32'd9; 
32'd962: dataIn2 = 32'd53; 
32'd963: dataIn2 = 32'd1; 
32'd964: dataIn2 = 32'd8; 
32'd965: dataIn2 = 32'd19; 
32'd966: dataIn2 = 32'd21; 
32'd967: dataIn2 = 32'd40; 
32'd968: dataIn2 = 32'd82; 
32'd969: dataIn2 = 32'd95; 
32'd970: dataIn2 = 32'd63; 
32'd971: dataIn2 = 32'd90; 
32'd972: dataIn2 = 32'd50; 
32'd973: dataIn2 = 32'd53; 
32'd974: dataIn2 = 32'd47; 
32'd975: dataIn2 = 32'd5; 
32'd976: dataIn2 = 32'd88; 
32'd977: dataIn2 = 32'd53; 
32'd978: dataIn2 = 32'd14; 
32'd979: dataIn2 = 32'd59; 
32'd980: dataIn2 = 32'd28; 
32'd981: dataIn2 = 32'd88; 
32'd982: dataIn2 = 32'd40; 
32'd983: dataIn2 = 32'd99; 
32'd984: dataIn2 = 32'd14; 
32'd985: dataIn2 = 32'd37; 
32'd986: dataIn2 = 32'd47; 
32'd987: dataIn2 = 32'd100; 
32'd988: dataIn2 = 32'd23; 
32'd989: dataIn2 = 32'd75; 
32'd990: dataIn2 = 32'd28; 
32'd991: dataIn2 = 32'd20; 
32'd992: dataIn2 = 32'd83; 
32'd993: dataIn2 = 32'd52; 
32'd994: dataIn2 = 32'd0; 
32'd995: dataIn2 = 32'd82; 
32'd996: dataIn2 = 32'd89; 
32'd997: dataIn2 = 32'd67; 
32'd998: dataIn2 = 32'd85; 
32'd999: dataIn2 = 32'd77; 
32'd1000: dataIn2 = 32'd81; 
32'd1001: dataIn2 = 32'd52; 
32'd1002: dataIn2 = 32'd8; 
32'd1003: dataIn2 = 32'd5; 
32'd1004: dataIn2 = 32'd28; 
32'd1005: dataIn2 = 32'd44; 
32'd1006: dataIn2 = 32'd10; 
32'd1007: dataIn2 = 32'd2; 
32'd1008: dataIn2 = 32'd31; 
32'd1009: dataIn2 = 32'd4; 
32'd1010: dataIn2 = 32'd34; 
32'd1011: dataIn2 = 32'd65; 
32'd1012: dataIn2 = 32'd73; 
32'd1013: dataIn2 = 32'd100; 
32'd1014: dataIn2 = 32'd98; 
32'd1015: dataIn2 = 32'd68; 
32'd1016: dataIn2 = 32'd93; 
32'd1017: dataIn2 = 32'd97; 
32'd1018: dataIn2 = 32'd100; 
32'd1019: dataIn2 = 32'd67; 
32'd1020: dataIn2 = 32'd77; 
32'd1021: dataIn2 = 32'd31; 
32'd1022: dataIn2 = 32'd9; 
32'd1023: dataIn2 = 32'd60; 
32'd1024: dataIn2 = 32'd78; 
32'd1025: dataIn2 = 32'd55; 
32'd1026: dataIn2 = 32'd3; 
32'd1027: dataIn2 = 32'd40; 
32'd1028: dataIn2 = 32'd68; 
32'd1029: dataIn2 = 32'd74; 
32'd1030: dataIn2 = 32'd94; 
32'd1031: dataIn2 = 32'd47; 
32'd1032: dataIn2 = 32'd77; 
32'd1033: dataIn2 = 32'd59; 
32'd1034: dataIn2 = 32'd20; 
32'd1035: dataIn2 = 32'd37; 
32'd1036: dataIn2 = 32'd89; 
32'd1037: dataIn2 = 32'd58; 
32'd1038: dataIn2 = 32'd41; 
32'd1039: dataIn2 = 32'd54; 
32'd1040: dataIn2 = 32'd12; 
32'd1041: dataIn2 = 32'd29; 
32'd1042: dataIn2 = 32'd26; 
32'd1043: dataIn2 = 32'd93; 
32'd1044: dataIn2 = 32'd20; 
32'd1045: dataIn2 = 32'd69; 
32'd1046: dataIn2 = 32'd14; 
32'd1047: dataIn2 = 32'd43; 
32'd1048: dataIn2 = 32'd51; 
32'd1049: dataIn2 = 32'd43; 
32'd1050: dataIn2 = 32'd14; 
32'd1051: dataIn2 = 32'd22; 
32'd1052: dataIn2 = 32'd4; 
32'd1053: dataIn2 = 32'd84; 
32'd1054: dataIn2 = 32'd100; 
32'd1055: dataIn2 = 32'd57; 
32'd1056: dataIn2 = 32'd68; 
32'd1057: dataIn2 = 32'd47; 
32'd1058: dataIn2 = 32'd87; 
32'd1059: dataIn2 = 32'd95; 
32'd1060: dataIn2 = 32'd20; 
32'd1061: dataIn2 = 32'd48; 
32'd1062: dataIn2 = 32'd43; 
32'd1063: dataIn2 = 32'd89; 
32'd1064: dataIn2 = 32'd95; 
32'd1065: dataIn2 = 32'd73; 
32'd1066: dataIn2 = 32'd19; 
32'd1067: dataIn2 = 32'd5; 
32'd1068: dataIn2 = 32'd18; 
32'd1069: dataIn2 = 32'd72; 
32'd1070: dataIn2 = 32'd88; 
32'd1071: dataIn2 = 32'd38; 
32'd1072: dataIn2 = 32'd86; 
32'd1073: dataIn2 = 32'd48; 
32'd1074: dataIn2 = 32'd66; 
32'd1075: dataIn2 = 32'd78; 
32'd1076: dataIn2 = 32'd9; 
32'd1077: dataIn2 = 32'd72; 
32'd1078: dataIn2 = 32'd43; 
32'd1079: dataIn2 = 32'd47; 
32'd1080: dataIn2 = 32'd4; 
32'd1081: dataIn2 = 32'd55; 
32'd1082: dataIn2 = 32'd74; 
32'd1083: dataIn2 = 32'd17; 
32'd1084: dataIn2 = 32'd4; 
32'd1085: dataIn2 = 32'd35; 
32'd1086: dataIn2 = 32'd11; 
32'd1087: dataIn2 = 32'd39; 
32'd1088: dataIn2 = 32'd22; 
32'd1089: dataIn2 = 32'd51; 
32'd1090: dataIn2 = 32'd69; 
32'd1091: dataIn2 = 32'd40; 
32'd1092: dataIn2 = 32'd60; 
32'd1093: dataIn2 = 32'd60; 
32'd1094: dataIn2 = 32'd5; 
32'd1095: dataIn2 = 32'd3; 
32'd1096: dataIn2 = 32'd99; 
32'd1097: dataIn2 = 32'd11; 
32'd1098: dataIn2 = 32'd85; 
32'd1099: dataIn2 = 32'd35; 
32'd1100: dataIn2 = 32'd89; 
32'd1101: dataIn2 = 32'd79; 
32'd1102: dataIn2 = 32'd93; 
32'd1103: dataIn2 = 32'd68; 
32'd1104: dataIn2 = 32'd3; 
32'd1105: dataIn2 = 32'd100; 
32'd1106: dataIn2 = 32'd9; 
32'd1107: dataIn2 = 32'd89; 
32'd1108: dataIn2 = 32'd87; 
32'd1109: dataIn2 = 32'd31; 
32'd1110: dataIn2 = 32'd88; 
32'd1111: dataIn2 = 32'd88; 
32'd1112: dataIn2 = 32'd64; 
32'd1113: dataIn2 = 32'd11; 
32'd1114: dataIn2 = 32'd86; 
32'd1115: dataIn2 = 32'd12; 
32'd1116: dataIn2 = 32'd100; 
32'd1117: dataIn2 = 32'd15; 
32'd1118: dataIn2 = 32'd32; 
32'd1119: dataIn2 = 32'd16; 
32'd1120: dataIn2 = 32'd59; 
32'd1121: dataIn2 = 32'd36; 
32'd1122: dataIn2 = 32'd64; 
32'd1123: dataIn2 = 32'd21; 
32'd1124: dataIn2 = 32'd8; 
32'd1125: dataIn2 = 32'd6; 
32'd1126: dataIn2 = 32'd70; 
32'd1127: dataIn2 = 32'd39; 
32'd1128: dataIn2 = 32'd88; 
32'd1129: dataIn2 = 32'd52; 
32'd1130: dataIn2 = 32'd10; 
32'd1131: dataIn2 = 32'd87; 
32'd1132: dataIn2 = 32'd61; 
32'd1133: dataIn2 = 32'd22; 
32'd1134: dataIn2 = 32'd37; 
32'd1135: dataIn2 = 32'd42; 
32'd1136: dataIn2 = 32'd97; 
32'd1137: dataIn2 = 32'd73; 
32'd1138: dataIn2 = 32'd58; 
32'd1139: dataIn2 = 32'd100; 
32'd1140: dataIn2 = 32'd39; 
32'd1141: dataIn2 = 32'd27; 
32'd1142: dataIn2 = 32'd85; 
32'd1143: dataIn2 = 32'd63; 
32'd1144: dataIn2 = 32'd44; 
32'd1145: dataIn2 = 32'd46; 
32'd1146: dataIn2 = 32'd5; 
32'd1147: dataIn2 = 32'd62; 
32'd1148: dataIn2 = 32'd50; 
32'd1149: dataIn2 = 32'd91; 
32'd1150: dataIn2 = 32'd97; 
32'd1151: dataIn2 = 32'd23; 
32'd1152: dataIn2 = 32'd10; 
32'd1153: dataIn2 = 32'd77; 
32'd1154: dataIn2 = 32'd93; 
32'd1155: dataIn2 = 32'd48; 
32'd1156: dataIn2 = 32'd39; 
32'd1157: dataIn2 = 32'd61; 
32'd1158: dataIn2 = 32'd21; 
32'd1159: dataIn2 = 32'd90; 
32'd1160: dataIn2 = 32'd60; 
32'd1161: dataIn2 = 32'd65; 
32'd1162: dataIn2 = 32'd63; 
32'd1163: dataIn2 = 32'd28; 
32'd1164: dataIn2 = 32'd38; 
32'd1165: dataIn2 = 32'd57; 
32'd1166: dataIn2 = 32'd28; 
32'd1167: dataIn2 = 32'd74; 
32'd1168: dataIn2 = 32'd20; 
32'd1169: dataIn2 = 32'd8; 
32'd1170: dataIn2 = 32'd6; 
32'd1171: dataIn2 = 32'd63; 
32'd1172: dataIn2 = 32'd76; 
32'd1173: dataIn2 = 32'd58; 
32'd1174: dataIn2 = 32'd25; 
32'd1175: dataIn2 = 32'd10; 
32'd1176: dataIn2 = 32'd33; 
32'd1177: dataIn2 = 32'd1; 
32'd1178: dataIn2 = 32'd11; 
32'd1179: dataIn2 = 32'd53; 
32'd1180: dataIn2 = 32'd80; 
32'd1181: dataIn2 = 32'd99; 
32'd1182: dataIn2 = 32'd89; 
32'd1183: dataIn2 = 32'd30; 
32'd1184: dataIn2 = 32'd60; 
32'd1185: dataIn2 = 32'd9; 
32'd1186: dataIn2 = 32'd90; 
32'd1187: dataIn2 = 32'd23; 
32'd1188: dataIn2 = 32'd13; 
32'd1189: dataIn2 = 32'd24; 
32'd1190: dataIn2 = 32'd22; 
32'd1191: dataIn2 = 32'd60; 
32'd1192: dataIn2 = 32'd96; 
32'd1193: dataIn2 = 32'd84; 
32'd1194: dataIn2 = 32'd77; 
32'd1195: dataIn2 = 32'd54; 
32'd1196: dataIn2 = 32'd22; 
32'd1197: dataIn2 = 32'd91; 
32'd1198: dataIn2 = 32'd91; 
32'd1199: dataIn2 = 32'd99; 
32'd1200: dataIn2 = 32'd80; 
32'd1201: dataIn2 = 32'd73; 
32'd1202: dataIn2 = 32'd69; 
32'd1203: dataIn2 = 32'd57; 
32'd1204: dataIn2 = 32'd39; 
32'd1205: dataIn2 = 32'd3; 
32'd1206: dataIn2 = 32'd73; 
32'd1207: dataIn2 = 32'd55; 
32'd1208: dataIn2 = 32'd27; 
32'd1209: dataIn2 = 32'd46; 
32'd1210: dataIn2 = 32'd42; 
32'd1211: dataIn2 = 32'd81; 
32'd1212: dataIn2 = 32'd16; 
32'd1213: dataIn2 = 32'd65; 
32'd1214: dataIn2 = 32'd91; 
32'd1215: dataIn2 = 32'd72; 
32'd1216: dataIn2 = 32'd80; 
32'd1217: dataIn2 = 32'd29; 
32'd1218: dataIn2 = 32'd86; 
32'd1219: dataIn2 = 32'd42; 
32'd1220: dataIn2 = 32'd71; 
32'd1221: dataIn2 = 32'd18; 
32'd1222: dataIn2 = 32'd31; 
32'd1223: dataIn2 = 32'd32; 
32'd1224: dataIn2 = 32'd45; 
32'd1225: dataIn2 = 32'd10; 
32'd1226: dataIn2 = 32'd22; 
32'd1227: dataIn2 = 32'd26; 
32'd1228: dataIn2 = 32'd61; 
32'd1229: dataIn2 = 32'd3; 
32'd1230: dataIn2 = 32'd52; 
32'd1231: dataIn2 = 32'd90; 
32'd1232: dataIn2 = 32'd69; 
32'd1233: dataIn2 = 32'd32; 
32'd1234: dataIn2 = 32'd16; 
32'd1235: dataIn2 = 32'd75; 
32'd1236: dataIn2 = 32'd76; 
32'd1237: dataIn2 = 32'd11; 
32'd1238: dataIn2 = 32'd54; 
32'd1239: dataIn2 = 32'd8; 
32'd1240: dataIn2 = 32'd36; 
32'd1241: dataIn2 = 32'd68; 
32'd1242: dataIn2 = 32'd81; 
32'd1243: dataIn2 = 32'd45; 
32'd1244: dataIn2 = 32'd60; 
32'd1245: dataIn2 = 32'd86; 
32'd1246: dataIn2 = 32'd68; 
32'd1247: dataIn2 = 32'd37; 
32'd1248: dataIn2 = 32'd63; 
32'd1249: dataIn2 = 32'd2; 
32'd1250: dataIn2 = 32'd47; 
32'd1251: dataIn2 = 32'd6; 
32'd1252: dataIn2 = 32'd44; 
32'd1253: dataIn2 = 32'd14; 
32'd1254: dataIn2 = 32'd7; 
32'd1255: dataIn2 = 32'd1; 
32'd1256: dataIn2 = 32'd9; 
32'd1257: dataIn2 = 32'd97; 
32'd1258: dataIn2 = 32'd83; 
32'd1259: dataIn2 = 32'd98; 
32'd1260: dataIn2 = 32'd33; 
32'd1261: dataIn2 = 32'd62; 
32'd1262: dataIn2 = 32'd94; 
32'd1263: dataIn2 = 32'd29; 
32'd1264: dataIn2 = 32'd1; 
32'd1265: dataIn2 = 32'd91; 
32'd1266: dataIn2 = 32'd94; 
32'd1267: dataIn2 = 32'd55; 
32'd1268: dataIn2 = 32'd84; 
32'd1269: dataIn2 = 32'd91; 
32'd1270: dataIn2 = 32'd90; 
32'd1271: dataIn2 = 32'd46; 
32'd1272: dataIn2 = 32'd93; 
32'd1273: dataIn2 = 32'd80; 
32'd1274: dataIn2 = 32'd74; 
32'd1275: dataIn2 = 32'd17; 
32'd1276: dataIn2 = 32'd13; 
32'd1277: dataIn2 = 32'd27; 
32'd1278: dataIn2 = 32'd86; 
32'd1279: dataIn2 = 32'd1; 
32'd1280: dataIn2 = 32'd8; 
32'd1281: dataIn2 = 32'd44; 
32'd1282: dataIn2 = 32'd42; 
32'd1283: dataIn2 = 32'd77; 
32'd1284: dataIn2 = 32'd53; 
32'd1285: dataIn2 = 32'd35; 
32'd1286: dataIn2 = 32'd33; 
32'd1287: dataIn2 = 32'd80; 
32'd1288: dataIn2 = 32'd46; 
32'd1289: dataIn2 = 32'd44; 
32'd1290: dataIn2 = 32'd81; 
32'd1291: dataIn2 = 32'd40; 
32'd1292: dataIn2 = 32'd74; 
32'd1293: dataIn2 = 32'd92; 
32'd1294: dataIn2 = 32'd77; 
32'd1295: dataIn2 = 32'd15; 
32'd1296: dataIn2 = 32'd100; 
32'd1297: dataIn2 = 32'd20; 
32'd1298: dataIn2 = 32'd84; 
32'd1299: dataIn2 = 32'd30; 
32'd1300: dataIn2 = 32'd33; 
32'd1301: dataIn2 = 32'd66; 
32'd1302: dataIn2 = 32'd62; 
32'd1303: dataIn2 = 32'd70; 
32'd1304: dataIn2 = 32'd100; 
32'd1305: dataIn2 = 32'd10; 
32'd1306: dataIn2 = 32'd30; 
32'd1307: dataIn2 = 32'd72; 
32'd1308: dataIn2 = 32'd24; 
32'd1309: dataIn2 = 32'd26; 
32'd1310: dataIn2 = 32'd8; 
32'd1311: dataIn2 = 32'd68; 
32'd1312: dataIn2 = 32'd7; 
32'd1313: dataIn2 = 32'd98; 
32'd1314: dataIn2 = 32'd76; 
32'd1315: dataIn2 = 32'd82; 
32'd1316: dataIn2 = 32'd23; 
32'd1317: dataIn2 = 32'd48; 
32'd1318: dataIn2 = 32'd12; 
32'd1319: dataIn2 = 32'd83; 
32'd1320: dataIn2 = 32'd50; 
32'd1321: dataIn2 = 32'd97; 
32'd1322: dataIn2 = 32'd66; 
32'd1323: dataIn2 = 32'd40; 
32'd1324: dataIn2 = 32'd13; 
32'd1325: dataIn2 = 32'd28; 
32'd1326: dataIn2 = 32'd76; 
32'd1327: dataIn2 = 32'd41; 
32'd1328: dataIn2 = 32'd29; 
32'd1329: dataIn2 = 32'd56; 
32'd1330: dataIn2 = 32'd74; 
32'd1331: dataIn2 = 32'd22; 
32'd1332: dataIn2 = 32'd46; 
32'd1333: dataIn2 = 32'd64; 
32'd1334: dataIn2 = 32'd10; 
32'd1335: dataIn2 = 32'd98; 
32'd1336: dataIn2 = 32'd81; 
32'd1337: dataIn2 = 32'd74; 
32'd1338: dataIn2 = 32'd13; 
32'd1339: dataIn2 = 32'd38; 
32'd1340: dataIn2 = 32'd25; 
32'd1341: dataIn2 = 32'd31; 
32'd1342: dataIn2 = 32'd8; 
32'd1343: dataIn2 = 32'd73; 
32'd1344: dataIn2 = 32'd83; 
32'd1345: dataIn2 = 32'd85; 
32'd1346: dataIn2 = 32'd99; 
32'd1347: dataIn2 = 32'd2; 
32'd1348: dataIn2 = 32'd8; 
32'd1349: dataIn2 = 32'd64; 
32'd1350: dataIn2 = 32'd37; 
32'd1351: dataIn2 = 32'd50; 
32'd1352: dataIn2 = 32'd26; 
32'd1353: dataIn2 = 32'd20; 
32'd1354: dataIn2 = 32'd59; 
32'd1355: dataIn2 = 32'd14; 
32'd1356: dataIn2 = 32'd9; 
32'd1357: dataIn2 = 32'd65; 
32'd1358: dataIn2 = 32'd94; 
32'd1359: dataIn2 = 32'd25; 
32'd1360: dataIn2 = 32'd23; 
32'd1361: dataIn2 = 32'd39; 
32'd1362: dataIn2 = 32'd2; 
32'd1363: dataIn2 = 32'd12; 
32'd1364: dataIn2 = 32'd17; 
32'd1365: dataIn2 = 32'd73; 
32'd1366: dataIn2 = 32'd86; 
32'd1367: dataIn2 = 32'd0; 
32'd1368: dataIn2 = 32'd7; 
32'd1369: dataIn2 = 32'd53; 
32'd1370: dataIn2 = 32'd30; 
32'd1371: dataIn2 = 32'd7; 
32'd1372: dataIn2 = 32'd73; 
32'd1373: dataIn2 = 32'd9; 
32'd1374: dataIn2 = 32'd97; 
32'd1375: dataIn2 = 32'd85; 
32'd1376: dataIn2 = 32'd58; 
32'd1377: dataIn2 = 32'd57; 
32'd1378: dataIn2 = 32'd78; 
32'd1379: dataIn2 = 32'd91; 
32'd1380: dataIn2 = 32'd71; 
32'd1381: dataIn2 = 32'd20; 
32'd1382: dataIn2 = 32'd69; 
32'd1383: dataIn2 = 32'd70; 
32'd1384: dataIn2 = 32'd79; 
32'd1385: dataIn2 = 32'd1; 
32'd1386: dataIn2 = 32'd100; 
32'd1387: dataIn2 = 32'd0; 
32'd1388: dataIn2 = 32'd14; 
32'd1389: dataIn2 = 32'd16; 
32'd1390: dataIn2 = 32'd78; 
32'd1391: dataIn2 = 32'd7; 
32'd1392: dataIn2 = 32'd22; 
32'd1393: dataIn2 = 32'd23; 
32'd1394: dataIn2 = 32'd73; 
32'd1395: dataIn2 = 32'd28; 
32'd1396: dataIn2 = 32'd92; 
32'd1397: dataIn2 = 32'd5; 
32'd1398: dataIn2 = 32'd72; 
32'd1399: dataIn2 = 32'd31; 
32'd1400: dataIn2 = 32'd72; 
32'd1401: dataIn2 = 32'd15; 
32'd1402: dataIn2 = 32'd94; 
32'd1403: dataIn2 = 32'd14; 
32'd1404: dataIn2 = 32'd19; 
32'd1405: dataIn2 = 32'd24; 
32'd1406: dataIn2 = 32'd60; 
32'd1407: dataIn2 = 32'd49; 
32'd1408: dataIn2 = 32'd25; 
32'd1409: dataIn2 = 32'd89; 
32'd1410: dataIn2 = 32'd16; 
32'd1411: dataIn2 = 32'd69; 
32'd1412: dataIn2 = 32'd44; 
32'd1413: dataIn2 = 32'd77; 
32'd1414: dataIn2 = 32'd98; 
32'd1415: dataIn2 = 32'd64; 
32'd1416: dataIn2 = 32'd52; 
32'd1417: dataIn2 = 32'd4; 
32'd1418: dataIn2 = 32'd54; 
32'd1419: dataIn2 = 32'd25; 
32'd1420: dataIn2 = 32'd72; 
32'd1421: dataIn2 = 32'd29; 
32'd1422: dataIn2 = 32'd87; 
32'd1423: dataIn2 = 32'd54; 
32'd1424: dataIn2 = 32'd8; 
32'd1425: dataIn2 = 32'd76; 
32'd1426: dataIn2 = 32'd71; 
32'd1427: dataIn2 = 32'd52; 
32'd1428: dataIn2 = 32'd62; 
32'd1429: dataIn2 = 32'd4; 
32'd1430: dataIn2 = 32'd22; 
32'd1431: dataIn2 = 32'd24; 
32'd1432: dataIn2 = 32'd74; 
32'd1433: dataIn2 = 32'd12; 
32'd1434: dataIn2 = 32'd6; 
32'd1435: dataIn2 = 32'd100; 
32'd1436: dataIn2 = 32'd35; 
32'd1437: dataIn2 = 32'd54; 
32'd1438: dataIn2 = 32'd1; 
32'd1439: dataIn2 = 32'd42; 
32'd1440: dataIn2 = 32'd22; 
32'd1441: dataIn2 = 32'd82; 
32'd1442: dataIn2 = 32'd26; 
32'd1443: dataIn2 = 32'd13; 
32'd1444: dataIn2 = 32'd79; 
32'd1445: dataIn2 = 32'd18; 
32'd1446: dataIn2 = 32'd54; 
32'd1447: dataIn2 = 32'd97; 
32'd1448: dataIn2 = 32'd77; 
32'd1449: dataIn2 = 32'd88; 
32'd1450: dataIn2 = 32'd90; 
32'd1451: dataIn2 = 32'd82; 
32'd1452: dataIn2 = 32'd65; 
32'd1453: dataIn2 = 32'd7; 
32'd1454: dataIn2 = 32'd88; 
32'd1455: dataIn2 = 32'd32; 
32'd1456: dataIn2 = 32'd48; 
32'd1457: dataIn2 = 32'd27; 
32'd1458: dataIn2 = 32'd43; 
32'd1459: dataIn2 = 32'd93; 
32'd1460: dataIn2 = 32'd31; 
32'd1461: dataIn2 = 32'd93; 
32'd1462: dataIn2 = 32'd7; 
32'd1463: dataIn2 = 32'd17; 
32'd1464: dataIn2 = 32'd20; 
32'd1465: dataIn2 = 32'd44; 
32'd1466: dataIn2 = 32'd38; 
32'd1467: dataIn2 = 32'd9; 
32'd1468: dataIn2 = 32'd81; 
32'd1469: dataIn2 = 32'd35; 
32'd1470: dataIn2 = 32'd87; 
32'd1471: dataIn2 = 32'd0; 
32'd1472: dataIn2 = 32'd30; 
32'd1473: dataIn2 = 32'd42; 
32'd1474: dataIn2 = 32'd57; 
32'd1475: dataIn2 = 32'd59; 
32'd1476: dataIn2 = 32'd78; 
32'd1477: dataIn2 = 32'd93; 
32'd1478: dataIn2 = 32'd39; 
32'd1479: dataIn2 = 32'd54; 
32'd1480: dataIn2 = 32'd5; 
32'd1481: dataIn2 = 32'd44; 
32'd1482: dataIn2 = 32'd95; 
32'd1483: dataIn2 = 32'd98; 
32'd1484: dataIn2 = 32'd76; 
32'd1485: dataIn2 = 32'd12; 
32'd1486: dataIn2 = 32'd77; 
32'd1487: dataIn2 = 32'd22; 
32'd1488: dataIn2 = 32'd18; 
32'd1489: dataIn2 = 32'd59; 
32'd1490: dataIn2 = 32'd46; 
32'd1491: dataIn2 = 32'd44; 
32'd1492: dataIn2 = 32'd14; 
32'd1493: dataIn2 = 32'd89; 
32'd1494: dataIn2 = 32'd15; 
32'd1495: dataIn2 = 32'd36; 
32'd1496: dataIn2 = 32'd99; 
32'd1497: dataIn2 = 32'd19; 
32'd1498: dataIn2 = 32'd51; 
32'd1499: dataIn2 = 32'd48; 
32'd1500: dataIn2 = 32'd81; 
32'd1501: dataIn2 = 32'd38; 
32'd1502: dataIn2 = 32'd19; 
32'd1503: dataIn2 = 32'd90; 
32'd1504: dataIn2 = 32'd15; 
32'd1505: dataIn2 = 32'd24; 
32'd1506: dataIn2 = 32'd90; 
32'd1507: dataIn2 = 32'd35; 
32'd1508: dataIn2 = 32'd61; 
32'd1509: dataIn2 = 32'd34; 
32'd1510: dataIn2 = 32'd47; 
32'd1511: dataIn2 = 32'd83; 
32'd1512: dataIn2 = 32'd15; 
32'd1513: dataIn2 = 32'd93; 
32'd1514: dataIn2 = 32'd41; 
32'd1515: dataIn2 = 32'd93; 
32'd1516: dataIn2 = 32'd20; 
32'd1517: dataIn2 = 32'd23; 
32'd1518: dataIn2 = 32'd46; 
32'd1519: dataIn2 = 32'd20; 
32'd1520: dataIn2 = 32'd99; 
32'd1521: dataIn2 = 32'd14; 
32'd1522: dataIn2 = 32'd27; 
32'd1523: dataIn2 = 32'd4; 
32'd1524: dataIn2 = 32'd74; 
32'd1525: dataIn2 = 32'd0; 
32'd1526: dataIn2 = 32'd75; 
32'd1527: dataIn2 = 32'd15; 
32'd1528: dataIn2 = 32'd21; 
32'd1529: dataIn2 = 32'd91; 
32'd1530: dataIn2 = 32'd42; 
32'd1531: dataIn2 = 32'd100; 
32'd1532: dataIn2 = 32'd11; 
32'd1533: dataIn2 = 32'd92; 
32'd1534: dataIn2 = 32'd63; 
32'd1535: dataIn2 = 32'd24; 
32'd1536: dataIn2 = 32'd82; 
32'd1537: dataIn2 = 32'd76; 
32'd1538: dataIn2 = 32'd80; 
32'd1539: dataIn2 = 32'd87; 
32'd1540: dataIn2 = 32'd99; 
32'd1541: dataIn2 = 32'd4; 
32'd1542: dataIn2 = 32'd88; 
32'd1543: dataIn2 = 32'd12; 
32'd1544: dataIn2 = 32'd78; 
32'd1545: dataIn2 = 32'd25; 
32'd1546: dataIn2 = 32'd88; 
32'd1547: dataIn2 = 32'd46; 
32'd1548: dataIn2 = 32'd15; 
32'd1549: dataIn2 = 32'd92; 
32'd1550: dataIn2 = 32'd12; 
32'd1551: dataIn2 = 32'd25; 
32'd1552: dataIn2 = 32'd42; 
32'd1553: dataIn2 = 32'd19; 
32'd1554: dataIn2 = 32'd13; 
32'd1555: dataIn2 = 32'd6; 
32'd1556: dataIn2 = 32'd97; 
32'd1557: dataIn2 = 32'd68; 
32'd1558: dataIn2 = 32'd1; 
32'd1559: dataIn2 = 32'd87; 
32'd1560: dataIn2 = 32'd27; 
32'd1561: dataIn2 = 32'd66; 
32'd1562: dataIn2 = 32'd92; 
32'd1563: dataIn2 = 32'd26; 
32'd1564: dataIn2 = 32'd88; 
32'd1565: dataIn2 = 32'd2; 
32'd1566: dataIn2 = 32'd6; 
32'd1567: dataIn2 = 32'd42; 
32'd1568: dataIn2 = 32'd43; 
32'd1569: dataIn2 = 32'd73; 
32'd1570: dataIn2 = 32'd54; 
32'd1571: dataIn2 = 32'd84; 
32'd1572: dataIn2 = 32'd79; 
32'd1573: dataIn2 = 32'd90; 
32'd1574: dataIn2 = 32'd62; 
32'd1575: dataIn2 = 32'd31; 
32'd1576: dataIn2 = 32'd40; 
32'd1577: dataIn2 = 32'd2; 
32'd1578: dataIn2 = 32'd88; 
32'd1579: dataIn2 = 32'd42; 
32'd1580: dataIn2 = 32'd42; 
32'd1581: dataIn2 = 32'd87; 
32'd1582: dataIn2 = 32'd6; 
32'd1583: dataIn2 = 32'd30; 
32'd1584: dataIn2 = 32'd55; 
32'd1585: dataIn2 = 32'd49; 
32'd1586: dataIn2 = 32'd48; 
32'd1587: dataIn2 = 32'd19; 
32'd1588: dataIn2 = 32'd9; 
32'd1589: dataIn2 = 32'd9; 
32'd1590: dataIn2 = 32'd49; 
32'd1591: dataIn2 = 32'd2; 
32'd1592: dataIn2 = 32'd51; 
32'd1593: dataIn2 = 32'd99; 
32'd1594: dataIn2 = 32'd49; 
32'd1595: dataIn2 = 32'd90; 
32'd1596: dataIn2 = 32'd70; 
32'd1597: dataIn2 = 32'd51; 
32'd1598: dataIn2 = 32'd0; 
32'd1599: dataIn2 = 32'd14; 
32'd1600: dataIn2 = 32'd15; 
32'd1601: dataIn2 = 32'd26; 
32'd1602: dataIn2 = 32'd53; 
32'd1603: dataIn2 = 32'd61; 
32'd1604: dataIn2 = 32'd13; 
32'd1605: dataIn2 = 32'd12; 
32'd1606: dataIn2 = 32'd23; 
32'd1607: dataIn2 = 32'd85; 
32'd1608: dataIn2 = 32'd12; 
32'd1609: dataIn2 = 32'd11; 
32'd1610: dataIn2 = 32'd15; 
32'd1611: dataIn2 = 32'd10; 
32'd1612: dataIn2 = 32'd52; 
32'd1613: dataIn2 = 32'd92; 
32'd1614: dataIn2 = 32'd55; 
32'd1615: dataIn2 = 32'd57; 
32'd1616: dataIn2 = 32'd94; 
32'd1617: dataIn2 = 32'd73; 
32'd1618: dataIn2 = 32'd62; 
32'd1619: dataIn2 = 32'd78; 
32'd1620: dataIn2 = 32'd66; 
32'd1621: dataIn2 = 32'd32; 
32'd1622: dataIn2 = 32'd84; 
32'd1623: dataIn2 = 32'd99; 
32'd1624: dataIn2 = 32'd84; 
32'd1625: dataIn2 = 32'd47; 
32'd1626: dataIn2 = 32'd61; 
32'd1627: dataIn2 = 32'd16; 
32'd1628: dataIn2 = 32'd81; 
32'd1629: dataIn2 = 32'd69; 
32'd1630: dataIn2 = 32'd37; 
32'd1631: dataIn2 = 32'd52; 
32'd1632: dataIn2 = 32'd60; 
32'd1633: dataIn2 = 32'd1; 
32'd1634: dataIn2 = 32'd48; 
32'd1635: dataIn2 = 32'd67; 
32'd1636: dataIn2 = 32'd39; 
32'd1637: dataIn2 = 32'd11; 
32'd1638: dataIn2 = 32'd39; 
32'd1639: dataIn2 = 32'd81; 
32'd1640: dataIn2 = 32'd53; 
32'd1641: dataIn2 = 32'd96; 
32'd1642: dataIn2 = 32'd28; 
32'd1643: dataIn2 = 32'd60; 
32'd1644: dataIn2 = 32'd55; 
32'd1645: dataIn2 = 32'd99; 
32'd1646: dataIn2 = 32'd32; 
32'd1647: dataIn2 = 32'd38; 
32'd1648: dataIn2 = 32'd59; 
32'd1649: dataIn2 = 32'd69; 
32'd1650: dataIn2 = 32'd81; 
32'd1651: dataIn2 = 32'd100; 
32'd1652: dataIn2 = 32'd50; 
32'd1653: dataIn2 = 32'd98; 
32'd1654: dataIn2 = 32'd60; 
32'd1655: dataIn2 = 32'd11; 
32'd1656: dataIn2 = 32'd1; 
32'd1657: dataIn2 = 32'd41; 
32'd1658: dataIn2 = 32'd49; 
32'd1659: dataIn2 = 32'd3; 
32'd1660: dataIn2 = 32'd54; 
32'd1661: dataIn2 = 32'd0; 
32'd1662: dataIn2 = 32'd7; 
32'd1663: dataIn2 = 32'd12; 
32'd1664: dataIn2 = 32'd35; 
32'd1665: dataIn2 = 32'd88; 
32'd1666: dataIn2 = 32'd44; 
32'd1667: dataIn2 = 32'd56; 
32'd1668: dataIn2 = 32'd71; 
32'd1669: dataIn2 = 32'd85; 
32'd1670: dataIn2 = 32'd62; 
32'd1671: dataIn2 = 32'd53; 
32'd1672: dataIn2 = 32'd5; 
32'd1673: dataIn2 = 32'd93; 
32'd1674: dataIn2 = 32'd35; 
32'd1675: dataIn2 = 32'd36; 
32'd1676: dataIn2 = 32'd48; 
32'd1677: dataIn2 = 32'd52; 
32'd1678: dataIn2 = 32'd58; 
32'd1679: dataIn2 = 32'd12; 
32'd1680: dataIn2 = 32'd77; 
32'd1681: dataIn2 = 32'd69; 
32'd1682: dataIn2 = 32'd8; 
32'd1683: dataIn2 = 32'd55; 
32'd1684: dataIn2 = 32'd70; 
32'd1685: dataIn2 = 32'd1; 
32'd1686: dataIn2 = 32'd22; 
32'd1687: dataIn2 = 32'd32; 
32'd1688: dataIn2 = 32'd89; 
32'd1689: dataIn2 = 32'd58; 
32'd1690: dataIn2 = 32'd47; 
32'd1691: dataIn2 = 32'd20; 
32'd1692: dataIn2 = 32'd25; 
32'd1693: dataIn2 = 32'd38; 
32'd1694: dataIn2 = 32'd1; 
32'd1695: dataIn2 = 32'd43; 
32'd1696: dataIn2 = 32'd43; 
32'd1697: dataIn2 = 32'd21; 
32'd1698: dataIn2 = 32'd4; 
32'd1699: dataIn2 = 32'd65; 
32'd1700: dataIn2 = 32'd20; 
32'd1701: dataIn2 = 32'd76; 
32'd1702: dataIn2 = 32'd51; 
32'd1703: dataIn2 = 32'd63; 
32'd1704: dataIn2 = 32'd100; 
32'd1705: dataIn2 = 32'd79; 
32'd1706: dataIn2 = 32'd22; 
32'd1707: dataIn2 = 32'd73; 
32'd1708: dataIn2 = 32'd81; 
32'd1709: dataIn2 = 32'd94; 
32'd1710: dataIn2 = 32'd1; 
32'd1711: dataIn2 = 32'd72; 
32'd1712: dataIn2 = 32'd63; 
32'd1713: dataIn2 = 32'd92; 
32'd1714: dataIn2 = 32'd98; 
32'd1715: dataIn2 = 32'd79; 
32'd1716: dataIn2 = 32'd25; 
32'd1717: dataIn2 = 32'd55; 
32'd1718: dataIn2 = 32'd90; 
32'd1719: dataIn2 = 32'd44; 
32'd1720: dataIn2 = 32'd50; 
32'd1721: dataIn2 = 32'd59; 
32'd1722: dataIn2 = 32'd100; 
32'd1723: dataIn2 = 32'd3; 
32'd1724: dataIn2 = 32'd18; 
32'd1725: dataIn2 = 32'd93; 
32'd1726: dataIn2 = 32'd65; 
32'd1727: dataIn2 = 32'd28; 
32'd1728: dataIn2 = 32'd7; 
32'd1729: dataIn2 = 32'd90; 
32'd1730: dataIn2 = 32'd68; 
32'd1731: dataIn2 = 32'd61; 
32'd1732: dataIn2 = 32'd99; 
32'd1733: dataIn2 = 32'd95; 
32'd1734: dataIn2 = 32'd97; 
32'd1735: dataIn2 = 32'd66; 
32'd1736: dataIn2 = 32'd63; 
32'd1737: dataIn2 = 32'd35; 
32'd1738: dataIn2 = 32'd69; 
32'd1739: dataIn2 = 32'd99; 
32'd1740: dataIn2 = 32'd61; 
32'd1741: dataIn2 = 32'd95; 
32'd1742: dataIn2 = 32'd60; 
32'd1743: dataIn2 = 32'd55; 
32'd1744: dataIn2 = 32'd77; 
32'd1745: dataIn2 = 32'd32; 
32'd1746: dataIn2 = 32'd73; 
32'd1747: dataIn2 = 32'd26; 
32'd1748: dataIn2 = 32'd37; 
32'd1749: dataIn2 = 32'd24; 
32'd1750: dataIn2 = 32'd36; 
32'd1751: dataIn2 = 32'd57; 
32'd1752: dataIn2 = 32'd46; 
32'd1753: dataIn2 = 32'd6; 
32'd1754: dataIn2 = 32'd25; 
32'd1755: dataIn2 = 32'd15; 
32'd1756: dataIn2 = 32'd30; 
32'd1757: dataIn2 = 32'd28; 
32'd1758: dataIn2 = 32'd33; 
32'd1759: dataIn2 = 32'd44; 
32'd1760: dataIn2 = 32'd7; 
32'd1761: dataIn2 = 32'd20; 
32'd1762: dataIn2 = 32'd13; 
32'd1763: dataIn2 = 32'd48; 
32'd1764: dataIn2 = 32'd92; 
32'd1765: dataIn2 = 32'd55; 
32'd1766: dataIn2 = 32'd22; 
32'd1767: dataIn2 = 32'd22; 
32'd1768: dataIn2 = 32'd87; 
32'd1769: dataIn2 = 32'd77; 
32'd1770: dataIn2 = 32'd67; 
32'd1771: dataIn2 = 32'd42; 
32'd1772: dataIn2 = 32'd62; 
32'd1773: dataIn2 = 32'd4; 
32'd1774: dataIn2 = 32'd22; 
32'd1775: dataIn2 = 32'd9; 
32'd1776: dataIn2 = 32'd100; 
32'd1777: dataIn2 = 32'd25; 
32'd1778: dataIn2 = 32'd16; 
32'd1779: dataIn2 = 32'd55; 
32'd1780: dataIn2 = 32'd53; 
32'd1781: dataIn2 = 32'd76; 
32'd1782: dataIn2 = 32'd13; 
32'd1783: dataIn2 = 32'd92; 
32'd1784: dataIn2 = 32'd6; 
32'd1785: dataIn2 = 32'd87; 
32'd1786: dataIn2 = 32'd94; 
32'd1787: dataIn2 = 32'd11; 
32'd1788: dataIn2 = 32'd22; 
32'd1789: dataIn2 = 32'd13; 
32'd1790: dataIn2 = 32'd40; 
32'd1791: dataIn2 = 32'd2; 
32'd1792: dataIn2 = 32'd89; 
32'd1793: dataIn2 = 32'd0; 
32'd1794: dataIn2 = 32'd1; 
32'd1795: dataIn2 = 32'd97; 
32'd1796: dataIn2 = 32'd89; 
32'd1797: dataIn2 = 32'd99; 
32'd1798: dataIn2 = 32'd94; 
32'd1799: dataIn2 = 32'd87; 
32'd1800: dataIn2 = 32'd18; 
32'd1801: dataIn2 = 32'd63; 
32'd1802: dataIn2 = 32'd11; 
32'd1803: dataIn2 = 32'd64; 
32'd1804: dataIn2 = 32'd53; 
32'd1805: dataIn2 = 32'd66; 
32'd1806: dataIn2 = 32'd29; 
32'd1807: dataIn2 = 32'd90; 
32'd1808: dataIn2 = 32'd1; 
32'd1809: dataIn2 = 32'd86; 
32'd1810: dataIn2 = 32'd84; 
32'd1811: dataIn2 = 32'd98; 
32'd1812: dataIn2 = 32'd30; 
32'd1813: dataIn2 = 32'd47; 
32'd1814: dataIn2 = 32'd44; 
32'd1815: dataIn2 = 32'd97; 
32'd1816: dataIn2 = 32'd40; 
32'd1817: dataIn2 = 32'd42; 
32'd1818: dataIn2 = 32'd24; 
32'd1819: dataIn2 = 32'd45; 
32'd1820: dataIn2 = 32'd37; 
32'd1821: dataIn2 = 32'd40; 
32'd1822: dataIn2 = 32'd77; 
32'd1823: dataIn2 = 32'd91; 
32'd1824: dataIn2 = 32'd59; 
32'd1825: dataIn2 = 32'd86; 
32'd1826: dataIn2 = 32'd41; 
32'd1827: dataIn2 = 32'd51; 
32'd1828: dataIn2 = 32'd98; 
32'd1829: dataIn2 = 32'd17; 
32'd1830: dataIn2 = 32'd6; 
32'd1831: dataIn2 = 32'd15; 
32'd1832: dataIn2 = 32'd67; 
32'd1833: dataIn2 = 32'd76; 
32'd1834: dataIn2 = 32'd52; 
32'd1835: dataIn2 = 32'd70; 
32'd1836: dataIn2 = 32'd1; 
32'd1837: dataIn2 = 32'd60; 
32'd1838: dataIn2 = 32'd4; 
32'd1839: dataIn2 = 32'd39; 
32'd1840: dataIn2 = 32'd28; 
32'd1841: dataIn2 = 32'd46; 
32'd1842: dataIn2 = 32'd34; 
32'd1843: dataIn2 = 32'd8; 
32'd1844: dataIn2 = 32'd52; 
32'd1845: dataIn2 = 32'd30; 
32'd1846: dataIn2 = 32'd37; 
32'd1847: dataIn2 = 32'd11; 
32'd1848: dataIn2 = 32'd97; 
32'd1849: dataIn2 = 32'd61; 
32'd1850: dataIn2 = 32'd84; 
32'd1851: dataIn2 = 32'd96; 
32'd1852: dataIn2 = 32'd91; 
32'd1853: dataIn2 = 32'd87; 
32'd1854: dataIn2 = 32'd11; 
32'd1855: dataIn2 = 32'd43; 
32'd1856: dataIn2 = 32'd88; 
32'd1857: dataIn2 = 32'd91; 
32'd1858: dataIn2 = 32'd72; 
32'd1859: dataIn2 = 32'd8; 
32'd1860: dataIn2 = 32'd15; 
32'd1861: dataIn2 = 32'd6; 
32'd1862: dataIn2 = 32'd71; 
32'd1863: dataIn2 = 32'd36; 
32'd1864: dataIn2 = 32'd51; 
32'd1865: dataIn2 = 32'd17; 
32'd1866: dataIn2 = 32'd91; 
32'd1867: dataIn2 = 32'd74; 
32'd1868: dataIn2 = 32'd71; 
32'd1869: dataIn2 = 32'd16; 
32'd1870: dataIn2 = 32'd9; 
32'd1871: dataIn2 = 32'd97; 
32'd1872: dataIn2 = 32'd98; 
32'd1873: dataIn2 = 32'd92; 
32'd1874: dataIn2 = 32'd19; 
32'd1875: dataIn2 = 32'd74; 
32'd1876: dataIn2 = 32'd72; 
32'd1877: dataIn2 = 32'd28; 
32'd1878: dataIn2 = 32'd70; 
32'd1879: dataIn2 = 32'd43; 
32'd1880: dataIn2 = 32'd13; 
32'd1881: dataIn2 = 32'd40; 
32'd1882: dataIn2 = 32'd24; 
32'd1883: dataIn2 = 32'd10; 
32'd1884: dataIn2 = 32'd97; 
32'd1885: dataIn2 = 32'd47; 
32'd1886: dataIn2 = 32'd93; 
32'd1887: dataIn2 = 32'd61; 
32'd1888: dataIn2 = 32'd31; 
32'd1889: dataIn2 = 32'd17; 
32'd1890: dataIn2 = 32'd48; 
32'd1891: dataIn2 = 32'd37; 
32'd1892: dataIn2 = 32'd13; 
32'd1893: dataIn2 = 32'd20; 
32'd1894: dataIn2 = 32'd1; 
32'd1895: dataIn2 = 32'd71; 
32'd1896: dataIn2 = 32'd36; 
32'd1897: dataIn2 = 32'd45; 
32'd1898: dataIn2 = 32'd4; 
32'd1899: dataIn2 = 32'd29; 
32'd1900: dataIn2 = 32'd67; 
32'd1901: dataIn2 = 32'd62; 
32'd1902: dataIn2 = 32'd46; 
32'd1903: dataIn2 = 32'd63; 
32'd1904: dataIn2 = 32'd16; 
32'd1905: dataIn2 = 32'd13; 
32'd1906: dataIn2 = 32'd62; 
32'd1907: dataIn2 = 32'd38; 
32'd1908: dataIn2 = 32'd17; 
32'd1909: dataIn2 = 32'd13; 
32'd1910: dataIn2 = 32'd4; 
32'd1911: dataIn2 = 32'd52; 
32'd1912: dataIn2 = 32'd4; 
32'd1913: dataIn2 = 32'd23; 
32'd1914: dataIn2 = 32'd84; 
32'd1915: dataIn2 = 32'd71; 
32'd1916: dataIn2 = 32'd77; 
32'd1917: dataIn2 = 32'd84; 
32'd1918: dataIn2 = 32'd80; 
32'd1919: dataIn2 = 32'd35; 
32'd1920: dataIn2 = 32'd45; 
32'd1921: dataIn2 = 32'd48; 
32'd1922: dataIn2 = 32'd66; 
32'd1923: dataIn2 = 32'd79; 
32'd1924: dataIn2 = 32'd38; 
32'd1925: dataIn2 = 32'd57; 
32'd1926: dataIn2 = 32'd66; 
32'd1927: dataIn2 = 32'd16; 
32'd1928: dataIn2 = 32'd28; 
32'd1929: dataIn2 = 32'd74; 
32'd1930: dataIn2 = 32'd53; 
32'd1931: dataIn2 = 32'd36; 
32'd1932: dataIn2 = 32'd39; 
32'd1933: dataIn2 = 32'd93; 
32'd1934: dataIn2 = 32'd26; 
32'd1935: dataIn2 = 32'd42; 
32'd1936: dataIn2 = 32'd82; 
32'd1937: dataIn2 = 32'd95; 
32'd1938: dataIn2 = 32'd17; 
32'd1939: dataIn2 = 32'd75; 
32'd1940: dataIn2 = 32'd68; 
32'd1941: dataIn2 = 32'd32; 
32'd1942: dataIn2 = 32'd72; 
32'd1943: dataIn2 = 32'd37; 
32'd1944: dataIn2 = 32'd76; 
32'd1945: dataIn2 = 32'd43; 
32'd1946: dataIn2 = 32'd63; 
32'd1947: dataIn2 = 32'd45; 
32'd1948: dataIn2 = 32'd75; 
32'd1949: dataIn2 = 32'd10; 
32'd1950: dataIn2 = 32'd49; 
32'd1951: dataIn2 = 32'd9; 
32'd1952: dataIn2 = 32'd71; 
32'd1953: dataIn2 = 32'd75; 
32'd1954: dataIn2 = 32'd18; 
32'd1955: dataIn2 = 32'd20; 
32'd1956: dataIn2 = 32'd53; 
32'd1957: dataIn2 = 32'd26; 
32'd1958: dataIn2 = 32'd87; 
32'd1959: dataIn2 = 32'd64; 
32'd1960: dataIn2 = 32'd74; 
32'd1961: dataIn2 = 32'd55; 
32'd1962: dataIn2 = 32'd8; 
32'd1963: dataIn2 = 32'd36; 
32'd1964: dataIn2 = 32'd96; 
32'd1965: dataIn2 = 32'd77; 
32'd1966: dataIn2 = 32'd30; 
32'd1967: dataIn2 = 32'd45; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_64_60.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
