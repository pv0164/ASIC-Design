//32x32 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 819 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd170 ; 
  wdata_col_base = 32'd9890 ; 
  row_base = 32'd107090 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #16560; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd107090: dataIn1 = 32'd0
; 
32'd107091: dataIn1 = 32'd22
; 
32'd107092: dataIn1 = 32'd49
; 
32'd107093: dataIn1 = 32'd75
; 
32'd107094: dataIn1 = 32'd98
; 
32'd107095: dataIn1 = 32'd120
; 
32'd107096: dataIn1 = 32'd143
; 
32'd107097: dataIn1 = 32'd166
; 
32'd107098: dataIn1 = 32'd185
; 
32'd107099: dataIn1 = 32'd211
; 
32'd107100: dataIn1 = 32'd236
; 
32'd107101: dataIn1 = 32'd263
; 
32'd107102: dataIn1 = 32'd289
; 
32'd107103: dataIn1 = 32'd314
; 
32'd107104: dataIn1 = 32'd340
; 
32'd107105: dataIn1 = 32'd362
; 
32'd107106: dataIn1 = 32'd388
; 
32'd107107: dataIn1 = 32'd413
; 
32'd107108: dataIn1 = 32'd439
; 
32'd107109: dataIn1 = 32'd464
; 
32'd107110: dataIn1 = 32'd489
; 
32'd107111: dataIn1 = 32'd514
; 
32'd107112: dataIn1 = 32'd536
; 
32'd107113: dataIn1 = 32'd559
; 
32'd107114: dataIn1 = 32'd585
; 
32'd107115: dataIn1 = 32'd606
; 
32'd107116: dataIn1 = 32'd631
; 
32'd107117: dataIn1 = 32'd658
; 
32'd107118: dataIn1 = 32'd680
; 
32'd107119: dataIn1 = 32'd707
; 
32'd107120: dataIn1 = 32'd728
; 
32'd107121: dataIn1 = 32'd752
; 
32'd107122: dataIn1 = 32'd780
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd9890: dataIn1 = 32'd0
; 
32'd9891: dataIn1 = 32'd22
; 
32'd9892: dataIn1 = 32'd49
; 
32'd9893: dataIn1 = 32'd75
; 
32'd9894: dataIn1 = 32'd98
; 
32'd9895: dataIn1 = 32'd120
; 
32'd9896: dataIn1 = 32'd143
; 
32'd9897: dataIn1 = 32'd166
; 
32'd9898: dataIn1 = 32'd185
; 
32'd9899: dataIn1 = 32'd211
; 
32'd9900: dataIn1 = 32'd236
; 
32'd9901: dataIn1 = 32'd263
; 
32'd9902: dataIn1 = 32'd289
; 
32'd9903: dataIn1 = 32'd314
; 
32'd9904: dataIn1 = 32'd340
; 
32'd9905: dataIn1 = 32'd362
; 
32'd9906: dataIn1 = 32'd388
; 
32'd9907: dataIn1 = 32'd413
; 
32'd9908: dataIn1 = 32'd439
; 
32'd9909: dataIn1 = 32'd464
; 
32'd9910: dataIn1 = 32'd489
; 
32'd9911: dataIn1 = 32'd514
; 
32'd9912: dataIn1 = 32'd536
; 
32'd9913: dataIn1 = 32'd559
; 
32'd9914: dataIn1 = 32'd585
; 
32'd9915: dataIn1 = 32'd606
; 
32'd9916: dataIn1 = 32'd631
; 
32'd9917: dataIn1 = 32'd658
; 
32'd9918: dataIn1 = 32'd680
; 
32'd9919: dataIn1 = 32'd707
; 
32'd9920: dataIn1 = 32'd728
; 
32'd9921: dataIn1 = 32'd752
; 
32'd9922: dataIn1 = 32'd780
; 
32'd9923: dataIn1 = 32'd0
; 
32'd9924: dataIn1 = 32'd1
; 
32'd9925: dataIn1 = 32'd2
; 
32'd9926: dataIn1 = 32'd3
; 
32'd9927: dataIn1 = 32'd4
; 
32'd9928: dataIn1 = 32'd5
; 
32'd9929: dataIn1 = 32'd6
; 
32'd9930: dataIn1 = 32'd7
; 
32'd9931: dataIn1 = 32'd10
; 
32'd9932: dataIn1 = 32'd11
; 
32'd9933: dataIn1 = 32'd12
; 
32'd9934: dataIn1 = 32'd16
; 
32'd9935: dataIn1 = 32'd18
; 
32'd9936: dataIn1 = 32'd19
; 
32'd9937: dataIn1 = 32'd21
; 
32'd9938: dataIn1 = 32'd23
; 
32'd9939: dataIn1 = 32'd25
; 
32'd9940: dataIn1 = 32'd26
; 
32'd9941: dataIn1 = 32'd28
; 
32'd9942: dataIn1 = 32'd29
; 
32'd9943: dataIn1 = 32'd30
; 
32'd9944: dataIn1 = 32'd31
; 
32'd9945: dataIn1 = 32'd0
; 
32'd9946: dataIn1 = 32'd1
; 
32'd9947: dataIn1 = 32'd2
; 
32'd9948: dataIn1 = 32'd3
; 
32'd9949: dataIn1 = 32'd5
; 
32'd9950: dataIn1 = 32'd6
; 
32'd9951: dataIn1 = 32'd8
; 
32'd9952: dataIn1 = 32'd9
; 
32'd9953: dataIn1 = 32'd10
; 
32'd9954: dataIn1 = 32'd11
; 
32'd9955: dataIn1 = 32'd12
; 
32'd9956: dataIn1 = 32'd13
; 
32'd9957: dataIn1 = 32'd14
; 
32'd9958: dataIn1 = 32'd15
; 
32'd9959: dataIn1 = 32'd16
; 
32'd9960: dataIn1 = 32'd20
; 
32'd9961: dataIn1 = 32'd21
; 
32'd9962: dataIn1 = 32'd22
; 
32'd9963: dataIn1 = 32'd23
; 
32'd9964: dataIn1 = 32'd24
; 
32'd9965: dataIn1 = 32'd25
; 
32'd9966: dataIn1 = 32'd26
; 
32'd9967: dataIn1 = 32'd27
; 
32'd9968: dataIn1 = 32'd28
; 
32'd9969: dataIn1 = 32'd29
; 
32'd9970: dataIn1 = 32'd30
; 
32'd9971: dataIn1 = 32'd31
; 
32'd9972: dataIn1 = 32'd0
; 
32'd9973: dataIn1 = 32'd3
; 
32'd9974: dataIn1 = 32'd4
; 
32'd9975: dataIn1 = 32'd5
; 
32'd9976: dataIn1 = 32'd7
; 
32'd9977: dataIn1 = 32'd8
; 
32'd9978: dataIn1 = 32'd9
; 
32'd9979: dataIn1 = 32'd10
; 
32'd9980: dataIn1 = 32'd12
; 
32'd9981: dataIn1 = 32'd13
; 
32'd9982: dataIn1 = 32'd15
; 
32'd9983: dataIn1 = 32'd16
; 
32'd9984: dataIn1 = 32'd17
; 
32'd9985: dataIn1 = 32'd18
; 
32'd9986: dataIn1 = 32'd19
; 
32'd9987: dataIn1 = 32'd20
; 
32'd9988: dataIn1 = 32'd21
; 
32'd9989: dataIn1 = 32'd22
; 
32'd9990: dataIn1 = 32'd23
; 
32'd9991: dataIn1 = 32'd24
; 
32'd9992: dataIn1 = 32'd25
; 
32'd9993: dataIn1 = 32'd26
; 
32'd9994: dataIn1 = 32'd27
; 
32'd9995: dataIn1 = 32'd28
; 
32'd9996: dataIn1 = 32'd30
; 
32'd9997: dataIn1 = 32'd31
; 
32'd9998: dataIn1 = 32'd0
; 
32'd9999: dataIn1 = 32'd2
; 
32'd10000: dataIn1 = 32'd4
; 
32'd10001: dataIn1 = 32'd5
; 
32'd10002: dataIn1 = 32'd7
; 
32'd10003: dataIn1 = 32'd10
; 
32'd10004: dataIn1 = 32'd12
; 
32'd10005: dataIn1 = 32'd13
; 
32'd10006: dataIn1 = 32'd14
; 
32'd10007: dataIn1 = 32'd15
; 
32'd10008: dataIn1 = 32'd18
; 
32'd10009: dataIn1 = 32'd19
; 
32'd10010: dataIn1 = 32'd20
; 
32'd10011: dataIn1 = 32'd21
; 
32'd10012: dataIn1 = 32'd22
; 
32'd10013: dataIn1 = 32'd23
; 
32'd10014: dataIn1 = 32'd24
; 
32'd10015: dataIn1 = 32'd25
; 
32'd10016: dataIn1 = 32'd26
; 
32'd10017: dataIn1 = 32'd28
; 
32'd10018: dataIn1 = 32'd29
; 
32'd10019: dataIn1 = 32'd30
; 
32'd10020: dataIn1 = 32'd31
; 
32'd10021: dataIn1 = 32'd1
; 
32'd10022: dataIn1 = 32'd3
; 
32'd10023: dataIn1 = 32'd6
; 
32'd10024: dataIn1 = 32'd7
; 
32'd10025: dataIn1 = 32'd10
; 
32'd10026: dataIn1 = 32'd11
; 
32'd10027: dataIn1 = 32'd12
; 
32'd10028: dataIn1 = 32'd13
; 
32'd10029: dataIn1 = 32'd14
; 
32'd10030: dataIn1 = 32'd15
; 
32'd10031: dataIn1 = 32'd16
; 
32'd10032: dataIn1 = 32'd18
; 
32'd10033: dataIn1 = 32'd19
; 
32'd10034: dataIn1 = 32'd20
; 
32'd10035: dataIn1 = 32'd22
; 
32'd10036: dataIn1 = 32'd23
; 
32'd10037: dataIn1 = 32'd24
; 
32'd10038: dataIn1 = 32'd25
; 
32'd10039: dataIn1 = 32'd26
; 
32'd10040: dataIn1 = 32'd28
; 
32'd10041: dataIn1 = 32'd29
; 
32'd10042: dataIn1 = 32'd30
; 
32'd10043: dataIn1 = 32'd0
; 
32'd10044: dataIn1 = 32'd1
; 
32'd10045: dataIn1 = 32'd3
; 
32'd10046: dataIn1 = 32'd4
; 
32'd10047: dataIn1 = 32'd5
; 
32'd10048: dataIn1 = 32'd6
; 
32'd10049: dataIn1 = 32'd8
; 
32'd10050: dataIn1 = 32'd9
; 
32'd10051: dataIn1 = 32'd10
; 
32'd10052: dataIn1 = 32'd12
; 
32'd10053: dataIn1 = 32'd13
; 
32'd10054: dataIn1 = 32'd14
; 
32'd10055: dataIn1 = 32'd16
; 
32'd10056: dataIn1 = 32'd18
; 
32'd10057: dataIn1 = 32'd19
; 
32'd10058: dataIn1 = 32'd20
; 
32'd10059: dataIn1 = 32'd21
; 
32'd10060: dataIn1 = 32'd23
; 
32'd10061: dataIn1 = 32'd24
; 
32'd10062: dataIn1 = 32'd25
; 
32'd10063: dataIn1 = 32'd26
; 
32'd10064: dataIn1 = 32'd28
; 
32'd10065: dataIn1 = 32'd30
; 
32'd10066: dataIn1 = 32'd0
; 
32'd10067: dataIn1 = 32'd5
; 
32'd10068: dataIn1 = 32'd7
; 
32'd10069: dataIn1 = 32'd8
; 
32'd10070: dataIn1 = 32'd9
; 
32'd10071: dataIn1 = 32'd10
; 
32'd10072: dataIn1 = 32'd12
; 
32'd10073: dataIn1 = 32'd13
; 
32'd10074: dataIn1 = 32'd14
; 
32'd10075: dataIn1 = 32'd15
; 
32'd10076: dataIn1 = 32'd16
; 
32'd10077: dataIn1 = 32'd17
; 
32'd10078: dataIn1 = 32'd19
; 
32'd10079: dataIn1 = 32'd20
; 
32'd10080: dataIn1 = 32'd21
; 
32'd10081: dataIn1 = 32'd22
; 
32'd10082: dataIn1 = 32'd23
; 
32'd10083: dataIn1 = 32'd24
; 
32'd10084: dataIn1 = 32'd26
; 
32'd10085: dataIn1 = 32'd27
; 
32'd10086: dataIn1 = 32'd28
; 
32'd10087: dataIn1 = 32'd29
; 
32'd10088: dataIn1 = 32'd31
; 
32'd10089: dataIn1 = 32'd1
; 
32'd10090: dataIn1 = 32'd2
; 
32'd10091: dataIn1 = 32'd4
; 
32'd10092: dataIn1 = 32'd7
; 
32'd10093: dataIn1 = 32'd8
; 
32'd10094: dataIn1 = 32'd9
; 
32'd10095: dataIn1 = 32'd10
; 
32'd10096: dataIn1 = 32'd12
; 
32'd10097: dataIn1 = 32'd14
; 
32'd10098: dataIn1 = 32'd17
; 
32'd10099: dataIn1 = 32'd18
; 
32'd10100: dataIn1 = 32'd19
; 
32'd10101: dataIn1 = 32'd20
; 
32'd10102: dataIn1 = 32'd21
; 
32'd10103: dataIn1 = 32'd23
; 
32'd10104: dataIn1 = 32'd24
; 
32'd10105: dataIn1 = 32'd25
; 
32'd10106: dataIn1 = 32'd29
; 
32'd10107: dataIn1 = 32'd30
; 
32'd10108: dataIn1 = 32'd0
; 
32'd10109: dataIn1 = 32'd3
; 
32'd10110: dataIn1 = 32'd5
; 
32'd10111: dataIn1 = 32'd6
; 
32'd10112: dataIn1 = 32'd7
; 
32'd10113: dataIn1 = 32'd8
; 
32'd10114: dataIn1 = 32'd9
; 
32'd10115: dataIn1 = 32'd10
; 
32'd10116: dataIn1 = 32'd11
; 
32'd10117: dataIn1 = 32'd12
; 
32'd10118: dataIn1 = 32'd14
; 
32'd10119: dataIn1 = 32'd15
; 
32'd10120: dataIn1 = 32'd16
; 
32'd10121: dataIn1 = 32'd17
; 
32'd10122: dataIn1 = 32'd18
; 
32'd10123: dataIn1 = 32'd19
; 
32'd10124: dataIn1 = 32'd20
; 
32'd10125: dataIn1 = 32'd21
; 
32'd10126: dataIn1 = 32'd22
; 
32'd10127: dataIn1 = 32'd23
; 
32'd10128: dataIn1 = 32'd24
; 
32'd10129: dataIn1 = 32'd25
; 
32'd10130: dataIn1 = 32'd26
; 
32'd10131: dataIn1 = 32'd27
; 
32'd10132: dataIn1 = 32'd30
; 
32'd10133: dataIn1 = 32'd31
; 
32'd10134: dataIn1 = 32'd0
; 
32'd10135: dataIn1 = 32'd1
; 
32'd10136: dataIn1 = 32'd3
; 
32'd10137: dataIn1 = 32'd4
; 
32'd10138: dataIn1 = 32'd7
; 
32'd10139: dataIn1 = 32'd8
; 
32'd10140: dataIn1 = 32'd9
; 
32'd10141: dataIn1 = 32'd10
; 
32'd10142: dataIn1 = 32'd11
; 
32'd10143: dataIn1 = 32'd13
; 
32'd10144: dataIn1 = 32'd14
; 
32'd10145: dataIn1 = 32'd15
; 
32'd10146: dataIn1 = 32'd16
; 
32'd10147: dataIn1 = 32'd18
; 
32'd10148: dataIn1 = 32'd19
; 
32'd10149: dataIn1 = 32'd20
; 
32'd10150: dataIn1 = 32'd21
; 
32'd10151: dataIn1 = 32'd22
; 
32'd10152: dataIn1 = 32'd24
; 
32'd10153: dataIn1 = 32'd25
; 
32'd10154: dataIn1 = 32'd26
; 
32'd10155: dataIn1 = 32'd27
; 
32'd10156: dataIn1 = 32'd28
; 
32'd10157: dataIn1 = 32'd29
; 
32'd10158: dataIn1 = 32'd30
; 
32'd10159: dataIn1 = 32'd0
; 
32'd10160: dataIn1 = 32'd1
; 
32'd10161: dataIn1 = 32'd2
; 
32'd10162: dataIn1 = 32'd3
; 
32'd10163: dataIn1 = 32'd4
; 
32'd10164: dataIn1 = 32'd5
; 
32'd10165: dataIn1 = 32'd6
; 
32'd10166: dataIn1 = 32'd7
; 
32'd10167: dataIn1 = 32'd8
; 
32'd10168: dataIn1 = 32'd10
; 
32'd10169: dataIn1 = 32'd11
; 
32'd10170: dataIn1 = 32'd12
; 
32'd10171: dataIn1 = 32'd13
; 
32'd10172: dataIn1 = 32'd14
; 
32'd10173: dataIn1 = 32'd15
; 
32'd10174: dataIn1 = 32'd16
; 
32'd10175: dataIn1 = 32'd17
; 
32'd10176: dataIn1 = 32'd18
; 
32'd10177: dataIn1 = 32'd19
; 
32'd10178: dataIn1 = 32'd21
; 
32'd10179: dataIn1 = 32'd22
; 
32'd10180: dataIn1 = 32'd23
; 
32'd10181: dataIn1 = 32'd25
; 
32'd10182: dataIn1 = 32'd27
; 
32'd10183: dataIn1 = 32'd28
; 
32'd10184: dataIn1 = 32'd29
; 
32'd10185: dataIn1 = 32'd31
; 
32'd10186: dataIn1 = 32'd0
; 
32'd10187: dataIn1 = 32'd1
; 
32'd10188: dataIn1 = 32'd2
; 
32'd10189: dataIn1 = 32'd3
; 
32'd10190: dataIn1 = 32'd4
; 
32'd10191: dataIn1 = 32'd6
; 
32'd10192: dataIn1 = 32'd7
; 
32'd10193: dataIn1 = 32'd8
; 
32'd10194: dataIn1 = 32'd10
; 
32'd10195: dataIn1 = 32'd11
; 
32'd10196: dataIn1 = 32'd12
; 
32'd10197: dataIn1 = 32'd13
; 
32'd10198: dataIn1 = 32'd17
; 
32'd10199: dataIn1 = 32'd18
; 
32'd10200: dataIn1 = 32'd19
; 
32'd10201: dataIn1 = 32'd20
; 
32'd10202: dataIn1 = 32'd21
; 
32'd10203: dataIn1 = 32'd22
; 
32'd10204: dataIn1 = 32'd23
; 
32'd10205: dataIn1 = 32'd24
; 
32'd10206: dataIn1 = 32'd25
; 
32'd10207: dataIn1 = 32'd26
; 
32'd10208: dataIn1 = 32'd27
; 
32'd10209: dataIn1 = 32'd28
; 
32'd10210: dataIn1 = 32'd30
; 
32'd10211: dataIn1 = 32'd31
; 
32'd10212: dataIn1 = 32'd0
; 
32'd10213: dataIn1 = 32'd2
; 
32'd10214: dataIn1 = 32'd3
; 
32'd10215: dataIn1 = 32'd4
; 
32'd10216: dataIn1 = 32'd5
; 
32'd10217: dataIn1 = 32'd6
; 
32'd10218: dataIn1 = 32'd7
; 
32'd10219: dataIn1 = 32'd8
; 
32'd10220: dataIn1 = 32'd9
; 
32'd10221: dataIn1 = 32'd12
; 
32'd10222: dataIn1 = 32'd13
; 
32'd10223: dataIn1 = 32'd14
; 
32'd10224: dataIn1 = 32'd16
; 
32'd10225: dataIn1 = 32'd18
; 
32'd10226: dataIn1 = 32'd19
; 
32'd10227: dataIn1 = 32'd21
; 
32'd10228: dataIn1 = 32'd22
; 
32'd10229: dataIn1 = 32'd23
; 
32'd10230: dataIn1 = 32'd24
; 
32'd10231: dataIn1 = 32'd25
; 
32'd10232: dataIn1 = 32'd27
; 
32'd10233: dataIn1 = 32'd28
; 
32'd10234: dataIn1 = 32'd29
; 
32'd10235: dataIn1 = 32'd30
; 
32'd10236: dataIn1 = 32'd31
; 
32'd10237: dataIn1 = 32'd0
; 
32'd10238: dataIn1 = 32'd1
; 
32'd10239: dataIn1 = 32'd2
; 
32'd10240: dataIn1 = 32'd3
; 
32'd10241: dataIn1 = 32'd4
; 
32'd10242: dataIn1 = 32'd5
; 
32'd10243: dataIn1 = 32'd6
; 
32'd10244: dataIn1 = 32'd7
; 
32'd10245: dataIn1 = 32'd9
; 
32'd10246: dataIn1 = 32'd10
; 
32'd10247: dataIn1 = 32'd11
; 
32'd10248: dataIn1 = 32'd13
; 
32'd10249: dataIn1 = 32'd14
; 
32'd10250: dataIn1 = 32'd18
; 
32'd10251: dataIn1 = 32'd19
; 
32'd10252: dataIn1 = 32'd20
; 
32'd10253: dataIn1 = 32'd21
; 
32'd10254: dataIn1 = 32'd22
; 
32'd10255: dataIn1 = 32'd23
; 
32'd10256: dataIn1 = 32'd24
; 
32'd10257: dataIn1 = 32'd25
; 
32'd10258: dataIn1 = 32'd26
; 
32'd10259: dataIn1 = 32'd27
; 
32'd10260: dataIn1 = 32'd28
; 
32'd10261: dataIn1 = 32'd29
; 
32'd10262: dataIn1 = 32'd30
; 
32'd10263: dataIn1 = 32'd0
; 
32'd10264: dataIn1 = 32'd1
; 
32'd10265: dataIn1 = 32'd4
; 
32'd10266: dataIn1 = 32'd5
; 
32'd10267: dataIn1 = 32'd7
; 
32'd10268: dataIn1 = 32'd8
; 
32'd10269: dataIn1 = 32'd9
; 
32'd10270: dataIn1 = 32'd10
; 
32'd10271: dataIn1 = 32'd11
; 
32'd10272: dataIn1 = 32'd12
; 
32'd10273: dataIn1 = 32'd13
; 
32'd10274: dataIn1 = 32'd14
; 
32'd10275: dataIn1 = 32'd15
; 
32'd10276: dataIn1 = 32'd17
; 
32'd10277: dataIn1 = 32'd19
; 
32'd10278: dataIn1 = 32'd20
; 
32'd10279: dataIn1 = 32'd21
; 
32'd10280: dataIn1 = 32'd23
; 
32'd10281: dataIn1 = 32'd26
; 
32'd10282: dataIn1 = 32'd27
; 
32'd10283: dataIn1 = 32'd29
; 
32'd10284: dataIn1 = 32'd30
; 
32'd10285: dataIn1 = 32'd0
; 
32'd10286: dataIn1 = 32'd1
; 
32'd10287: dataIn1 = 32'd3
; 
32'd10288: dataIn1 = 32'd4
; 
32'd10289: dataIn1 = 32'd5
; 
32'd10290: dataIn1 = 32'd6
; 
32'd10291: dataIn1 = 32'd8
; 
32'd10292: dataIn1 = 32'd9
; 
32'd10293: dataIn1 = 32'd10
; 
32'd10294: dataIn1 = 32'd12
; 
32'd10295: dataIn1 = 32'd13
; 
32'd10296: dataIn1 = 32'd14
; 
32'd10297: dataIn1 = 32'd15
; 
32'd10298: dataIn1 = 32'd17
; 
32'd10299: dataIn1 = 32'd19
; 
32'd10300: dataIn1 = 32'd20
; 
32'd10301: dataIn1 = 32'd21
; 
32'd10302: dataIn1 = 32'd22
; 
32'd10303: dataIn1 = 32'd23
; 
32'd10304: dataIn1 = 32'd24
; 
32'd10305: dataIn1 = 32'd25
; 
32'd10306: dataIn1 = 32'd27
; 
32'd10307: dataIn1 = 32'd28
; 
32'd10308: dataIn1 = 32'd29
; 
32'd10309: dataIn1 = 32'd30
; 
32'd10310: dataIn1 = 32'd31
; 
32'd10311: dataIn1 = 32'd0
; 
32'd10312: dataIn1 = 32'd1
; 
32'd10313: dataIn1 = 32'd2
; 
32'd10314: dataIn1 = 32'd3
; 
32'd10315: dataIn1 = 32'd4
; 
32'd10316: dataIn1 = 32'd6
; 
32'd10317: dataIn1 = 32'd7
; 
32'd10318: dataIn1 = 32'd10
; 
32'd10319: dataIn1 = 32'd11
; 
32'd10320: dataIn1 = 32'd12
; 
32'd10321: dataIn1 = 32'd14
; 
32'd10322: dataIn1 = 32'd15
; 
32'd10323: dataIn1 = 32'd16
; 
32'd10324: dataIn1 = 32'd18
; 
32'd10325: dataIn1 = 32'd19
; 
32'd10326: dataIn1 = 32'd20
; 
32'd10327: dataIn1 = 32'd21
; 
32'd10328: dataIn1 = 32'd22
; 
32'd10329: dataIn1 = 32'd23
; 
32'd10330: dataIn1 = 32'd25
; 
32'd10331: dataIn1 = 32'd26
; 
32'd10332: dataIn1 = 32'd27
; 
32'd10333: dataIn1 = 32'd28
; 
32'd10334: dataIn1 = 32'd29
; 
32'd10335: dataIn1 = 32'd31
; 
32'd10336: dataIn1 = 32'd0
; 
32'd10337: dataIn1 = 32'd1
; 
32'd10338: dataIn1 = 32'd3
; 
32'd10339: dataIn1 = 32'd4
; 
32'd10340: dataIn1 = 32'd5
; 
32'd10341: dataIn1 = 32'd6
; 
32'd10342: dataIn1 = 32'd7
; 
32'd10343: dataIn1 = 32'd9
; 
32'd10344: dataIn1 = 32'd10
; 
32'd10345: dataIn1 = 32'd11
; 
32'd10346: dataIn1 = 32'd12
; 
32'd10347: dataIn1 = 32'd13
; 
32'd10348: dataIn1 = 32'd14
; 
32'd10349: dataIn1 = 32'd16
; 
32'd10350: dataIn1 = 32'd17
; 
32'd10351: dataIn1 = 32'd19
; 
32'd10352: dataIn1 = 32'd20
; 
32'd10353: dataIn1 = 32'd22
; 
32'd10354: dataIn1 = 32'd23
; 
32'd10355: dataIn1 = 32'd25
; 
32'd10356: dataIn1 = 32'd26
; 
32'd10357: dataIn1 = 32'd27
; 
32'd10358: dataIn1 = 32'd28
; 
32'd10359: dataIn1 = 32'd29
; 
32'd10360: dataIn1 = 32'd30
; 
32'd10361: dataIn1 = 32'd31
; 
32'd10362: dataIn1 = 32'd0
; 
32'd10363: dataIn1 = 32'd2
; 
32'd10364: dataIn1 = 32'd4
; 
32'd10365: dataIn1 = 32'd5
; 
32'd10366: dataIn1 = 32'd6
; 
32'd10367: dataIn1 = 32'd8
; 
32'd10368: dataIn1 = 32'd9
; 
32'd10369: dataIn1 = 32'd11
; 
32'd10370: dataIn1 = 32'd13
; 
32'd10371: dataIn1 = 32'd14
; 
32'd10372: dataIn1 = 32'd15
; 
32'd10373: dataIn1 = 32'd16
; 
32'd10374: dataIn1 = 32'd18
; 
32'd10375: dataIn1 = 32'd19
; 
32'd10376: dataIn1 = 32'd20
; 
32'd10377: dataIn1 = 32'd21
; 
32'd10378: dataIn1 = 32'd22
; 
32'd10379: dataIn1 = 32'd23
; 
32'd10380: dataIn1 = 32'd24
; 
32'd10381: dataIn1 = 32'd25
; 
32'd10382: dataIn1 = 32'd27
; 
32'd10383: dataIn1 = 32'd28
; 
32'd10384: dataIn1 = 32'd29
; 
32'd10385: dataIn1 = 32'd30
; 
32'd10386: dataIn1 = 32'd31
; 
32'd10387: dataIn1 = 32'd0
; 
32'd10388: dataIn1 = 32'd1
; 
32'd10389: dataIn1 = 32'd2
; 
32'd10390: dataIn1 = 32'd3
; 
32'd10391: dataIn1 = 32'd5
; 
32'd10392: dataIn1 = 32'd7
; 
32'd10393: dataIn1 = 32'd8
; 
32'd10394: dataIn1 = 32'd9
; 
32'd10395: dataIn1 = 32'd10
; 
32'd10396: dataIn1 = 32'd12
; 
32'd10397: dataIn1 = 32'd13
; 
32'd10398: dataIn1 = 32'd14
; 
32'd10399: dataIn1 = 32'd15
; 
32'd10400: dataIn1 = 32'd16
; 
32'd10401: dataIn1 = 32'd17
; 
32'd10402: dataIn1 = 32'd18
; 
32'd10403: dataIn1 = 32'd19
; 
32'd10404: dataIn1 = 32'd21
; 
32'd10405: dataIn1 = 32'd23
; 
32'd10406: dataIn1 = 32'd24
; 
32'd10407: dataIn1 = 32'd25
; 
32'd10408: dataIn1 = 32'd26
; 
32'd10409: dataIn1 = 32'd27
; 
32'd10410: dataIn1 = 32'd29
; 
32'd10411: dataIn1 = 32'd31
; 
32'd10412: dataIn1 = 32'd0
; 
32'd10413: dataIn1 = 32'd1
; 
32'd10414: dataIn1 = 32'd2
; 
32'd10415: dataIn1 = 32'd3
; 
32'd10416: dataIn1 = 32'd5
; 
32'd10417: dataIn1 = 32'd6
; 
32'd10418: dataIn1 = 32'd8
; 
32'd10419: dataIn1 = 32'd9
; 
32'd10420: dataIn1 = 32'd10
; 
32'd10421: dataIn1 = 32'd11
; 
32'd10422: dataIn1 = 32'd12
; 
32'd10423: dataIn1 = 32'd13
; 
32'd10424: dataIn1 = 32'd14
; 
32'd10425: dataIn1 = 32'd15
; 
32'd10426: dataIn1 = 32'd16
; 
32'd10427: dataIn1 = 32'd17
; 
32'd10428: dataIn1 = 32'd18
; 
32'd10429: dataIn1 = 32'd19
; 
32'd10430: dataIn1 = 32'd20
; 
32'd10431: dataIn1 = 32'd21
; 
32'd10432: dataIn1 = 32'd22
; 
32'd10433: dataIn1 = 32'd23
; 
32'd10434: dataIn1 = 32'd26
; 
32'd10435: dataIn1 = 32'd28
; 
32'd10436: dataIn1 = 32'd29
; 
32'd10437: dataIn1 = 32'd0
; 
32'd10438: dataIn1 = 32'd2
; 
32'd10439: dataIn1 = 32'd4
; 
32'd10440: dataIn1 = 32'd5
; 
32'd10441: dataIn1 = 32'd9
; 
32'd10442: dataIn1 = 32'd11
; 
32'd10443: dataIn1 = 32'd12
; 
32'd10444: dataIn1 = 32'd13
; 
32'd10445: dataIn1 = 32'd14
; 
32'd10446: dataIn1 = 32'd15
; 
32'd10447: dataIn1 = 32'd16
; 
32'd10448: dataIn1 = 32'd17
; 
32'd10449: dataIn1 = 32'd18
; 
32'd10450: dataIn1 = 32'd19
; 
32'd10451: dataIn1 = 32'd20
; 
32'd10452: dataIn1 = 32'd21
; 
32'd10453: dataIn1 = 32'd23
; 
32'd10454: dataIn1 = 32'd24
; 
32'd10455: dataIn1 = 32'd25
; 
32'd10456: dataIn1 = 32'd27
; 
32'd10457: dataIn1 = 32'd28
; 
32'd10458: dataIn1 = 32'd29
; 
32'd10459: dataIn1 = 32'd0
; 
32'd10460: dataIn1 = 32'd1
; 
32'd10461: dataIn1 = 32'd2
; 
32'd10462: dataIn1 = 32'd5
; 
32'd10463: dataIn1 = 32'd6
; 
32'd10464: dataIn1 = 32'd7
; 
32'd10465: dataIn1 = 32'd8
; 
32'd10466: dataIn1 = 32'd9
; 
32'd10467: dataIn1 = 32'd10
; 
32'd10468: dataIn1 = 32'd11
; 
32'd10469: dataIn1 = 32'd13
; 
32'd10470: dataIn1 = 32'd15
; 
32'd10471: dataIn1 = 32'd16
; 
32'd10472: dataIn1 = 32'd17
; 
32'd10473: dataIn1 = 32'd18
; 
32'd10474: dataIn1 = 32'd20
; 
32'd10475: dataIn1 = 32'd21
; 
32'd10476: dataIn1 = 32'd23
; 
32'd10477: dataIn1 = 32'd24
; 
32'd10478: dataIn1 = 32'd26
; 
32'd10479: dataIn1 = 32'd27
; 
32'd10480: dataIn1 = 32'd28
; 
32'd10481: dataIn1 = 32'd31
; 
32'd10482: dataIn1 = 32'd0
; 
32'd10483: dataIn1 = 32'd1
; 
32'd10484: dataIn1 = 32'd2
; 
32'd10485: dataIn1 = 32'd3
; 
32'd10486: dataIn1 = 32'd4
; 
32'd10487: dataIn1 = 32'd5
; 
32'd10488: dataIn1 = 32'd6
; 
32'd10489: dataIn1 = 32'd7
; 
32'd10490: dataIn1 = 32'd8
; 
32'd10491: dataIn1 = 32'd9
; 
32'd10492: dataIn1 = 32'd10
; 
32'd10493: dataIn1 = 32'd11
; 
32'd10494: dataIn1 = 32'd12
; 
32'd10495: dataIn1 = 32'd15
; 
32'd10496: dataIn1 = 32'd16
; 
32'd10497: dataIn1 = 32'd17
; 
32'd10498: dataIn1 = 32'd18
; 
32'd10499: dataIn1 = 32'd21
; 
32'd10500: dataIn1 = 32'd22
; 
32'd10501: dataIn1 = 32'd23
; 
32'd10502: dataIn1 = 32'd24
; 
32'd10503: dataIn1 = 32'd25
; 
32'd10504: dataIn1 = 32'd27
; 
32'd10505: dataIn1 = 32'd28
; 
32'd10506: dataIn1 = 32'd30
; 
32'd10507: dataIn1 = 32'd31
; 
32'd10508: dataIn1 = 32'd0
; 
32'd10509: dataIn1 = 32'd1
; 
32'd10510: dataIn1 = 32'd2
; 
32'd10511: dataIn1 = 32'd4
; 
32'd10512: dataIn1 = 32'd6
; 
32'd10513: dataIn1 = 32'd7
; 
32'd10514: dataIn1 = 32'd8
; 
32'd10515: dataIn1 = 32'd9
; 
32'd10516: dataIn1 = 32'd12
; 
32'd10517: dataIn1 = 32'd14
; 
32'd10518: dataIn1 = 32'd15
; 
32'd10519: dataIn1 = 32'd17
; 
32'd10520: dataIn1 = 32'd19
; 
32'd10521: dataIn1 = 32'd21
; 
32'd10522: dataIn1 = 32'd22
; 
32'd10523: dataIn1 = 32'd23
; 
32'd10524: dataIn1 = 32'd26
; 
32'd10525: dataIn1 = 32'd28
; 
32'd10526: dataIn1 = 32'd29
; 
32'd10527: dataIn1 = 32'd30
; 
32'd10528: dataIn1 = 32'd31
; 
32'd10529: dataIn1 = 32'd0
; 
32'd10530: dataIn1 = 32'd4
; 
32'd10531: dataIn1 = 32'd5
; 
32'd10532: dataIn1 = 32'd6
; 
32'd10533: dataIn1 = 32'd8
; 
32'd10534: dataIn1 = 32'd9
; 
32'd10535: dataIn1 = 32'd11
; 
32'd10536: dataIn1 = 32'd13
; 
32'd10537: dataIn1 = 32'd14
; 
32'd10538: dataIn1 = 32'd15
; 
32'd10539: dataIn1 = 32'd16
; 
32'd10540: dataIn1 = 32'd17
; 
32'd10541: dataIn1 = 32'd19
; 
32'd10542: dataIn1 = 32'd20
; 
32'd10543: dataIn1 = 32'd21
; 
32'd10544: dataIn1 = 32'd22
; 
32'd10545: dataIn1 = 32'd23
; 
32'd10546: dataIn1 = 32'd24
; 
32'd10547: dataIn1 = 32'd25
; 
32'd10548: dataIn1 = 32'd26
; 
32'd10549: dataIn1 = 32'd27
; 
32'd10550: dataIn1 = 32'd28
; 
32'd10551: dataIn1 = 32'd29
; 
32'd10552: dataIn1 = 32'd30
; 
32'd10553: dataIn1 = 32'd31
; 
32'd10554: dataIn1 = 32'd0
; 
32'd10555: dataIn1 = 32'd1
; 
32'd10556: dataIn1 = 32'd2
; 
32'd10557: dataIn1 = 32'd3
; 
32'd10558: dataIn1 = 32'd4
; 
32'd10559: dataIn1 = 32'd5
; 
32'd10560: dataIn1 = 32'd6
; 
32'd10561: dataIn1 = 32'd7
; 
32'd10562: dataIn1 = 32'd8
; 
32'd10563: dataIn1 = 32'd10
; 
32'd10564: dataIn1 = 32'd11
; 
32'd10565: dataIn1 = 32'd12
; 
32'd10566: dataIn1 = 32'd13
; 
32'd10567: dataIn1 = 32'd14
; 
32'd10568: dataIn1 = 32'd15
; 
32'd10569: dataIn1 = 32'd16
; 
32'd10570: dataIn1 = 32'd17
; 
32'd10571: dataIn1 = 32'd18
; 
32'd10572: dataIn1 = 32'd19
; 
32'd10573: dataIn1 = 32'd20
; 
32'd10574: dataIn1 = 32'd21
; 
32'd10575: dataIn1 = 32'd22
; 
32'd10576: dataIn1 = 32'd27
; 
32'd10577: dataIn1 = 32'd28
; 
32'd10578: dataIn1 = 32'd29
; 
32'd10579: dataIn1 = 32'd30
; 
32'd10580: dataIn1 = 32'd31
; 
32'd10581: dataIn1 = 32'd2
; 
32'd10582: dataIn1 = 32'd3
; 
32'd10583: dataIn1 = 32'd5
; 
32'd10584: dataIn1 = 32'd6
; 
32'd10585: dataIn1 = 32'd7
; 
32'd10586: dataIn1 = 32'd9
; 
32'd10587: dataIn1 = 32'd10
; 
32'd10588: dataIn1 = 32'd12
; 
32'd10589: dataIn1 = 32'd13
; 
32'd10590: dataIn1 = 32'd18
; 
32'd10591: dataIn1 = 32'd19
; 
32'd10592: dataIn1 = 32'd20
; 
32'd10593: dataIn1 = 32'd21
; 
32'd10594: dataIn1 = 32'd22
; 
32'd10595: dataIn1 = 32'd23
; 
32'd10596: dataIn1 = 32'd24
; 
32'd10597: dataIn1 = 32'd25
; 
32'd10598: dataIn1 = 32'd26
; 
32'd10599: dataIn1 = 32'd27
; 
32'd10600: dataIn1 = 32'd29
; 
32'd10601: dataIn1 = 32'd30
; 
32'd10602: dataIn1 = 32'd31
; 
32'd10603: dataIn1 = 32'd0
; 
32'd10604: dataIn1 = 32'd1
; 
32'd10605: dataIn1 = 32'd2
; 
32'd10606: dataIn1 = 32'd3
; 
32'd10607: dataIn1 = 32'd4
; 
32'd10608: dataIn1 = 32'd5
; 
32'd10609: dataIn1 = 32'd6
; 
32'd10610: dataIn1 = 32'd7
; 
32'd10611: dataIn1 = 32'd8
; 
32'd10612: dataIn1 = 32'd9
; 
32'd10613: dataIn1 = 32'd10
; 
32'd10614: dataIn1 = 32'd11
; 
32'd10615: dataIn1 = 32'd12
; 
32'd10616: dataIn1 = 32'd13
; 
32'd10617: dataIn1 = 32'd14
; 
32'd10618: dataIn1 = 32'd15
; 
32'd10619: dataIn1 = 32'd17
; 
32'd10620: dataIn1 = 32'd19
; 
32'd10621: dataIn1 = 32'd20
; 
32'd10622: dataIn1 = 32'd21
; 
32'd10623: dataIn1 = 32'd22
; 
32'd10624: dataIn1 = 32'd23
; 
32'd10625: dataIn1 = 32'd24
; 
32'd10626: dataIn1 = 32'd25
; 
32'd10627: dataIn1 = 32'd26
; 
32'd10628: dataIn1 = 32'd27
; 
32'd10629: dataIn1 = 32'd28
; 
32'd10630: dataIn1 = 32'd0
; 
32'd10631: dataIn1 = 32'd2
; 
32'd10632: dataIn1 = 32'd3
; 
32'd10633: dataIn1 = 32'd5
; 
32'd10634: dataIn1 = 32'd10
; 
32'd10635: dataIn1 = 32'd11
; 
32'd10636: dataIn1 = 32'd12
; 
32'd10637: dataIn1 = 32'd13
; 
32'd10638: dataIn1 = 32'd14
; 
32'd10639: dataIn1 = 32'd15
; 
32'd10640: dataIn1 = 32'd17
; 
32'd10641: dataIn1 = 32'd18
; 
32'd10642: dataIn1 = 32'd19
; 
32'd10643: dataIn1 = 32'd20
; 
32'd10644: dataIn1 = 32'd22
; 
32'd10645: dataIn1 = 32'd23
; 
32'd10646: dataIn1 = 32'd24
; 
32'd10647: dataIn1 = 32'd25
; 
32'd10648: dataIn1 = 32'd29
; 
32'd10649: dataIn1 = 32'd30
; 
32'd10650: dataIn1 = 32'd31
; 
32'd10651: dataIn1 = 32'd0
; 
32'd10652: dataIn1 = 32'd1
; 
32'd10653: dataIn1 = 32'd2
; 
32'd10654: dataIn1 = 32'd3
; 
32'd10655: dataIn1 = 32'd4
; 
32'd10656: dataIn1 = 32'd5
; 
32'd10657: dataIn1 = 32'd6
; 
32'd10658: dataIn1 = 32'd8
; 
32'd10659: dataIn1 = 32'd9
; 
32'd10660: dataIn1 = 32'd11
; 
32'd10661: dataIn1 = 32'd12
; 
32'd10662: dataIn1 = 32'd13
; 
32'd10663: dataIn1 = 32'd14
; 
32'd10664: dataIn1 = 32'd16
; 
32'd10665: dataIn1 = 32'd17
; 
32'd10666: dataIn1 = 32'd18
; 
32'd10667: dataIn1 = 32'd19
; 
32'd10668: dataIn1 = 32'd20
; 
32'd10669: dataIn1 = 32'd21
; 
32'd10670: dataIn1 = 32'd22
; 
32'd10671: dataIn1 = 32'd25
; 
32'd10672: dataIn1 = 32'd26
; 
32'd10673: dataIn1 = 32'd28
; 
32'd10674: dataIn1 = 32'd30
; 
32'd10675: dataIn1 = 32'd0
; 
32'd10676: dataIn1 = 32'd2
; 
32'd10677: dataIn1 = 32'd3
; 
32'd10678: dataIn1 = 32'd4
; 
32'd10679: dataIn1 = 32'd5
; 
32'd10680: dataIn1 = 32'd6
; 
32'd10681: dataIn1 = 32'd7
; 
32'd10682: dataIn1 = 32'd8
; 
32'd10683: dataIn1 = 32'd9
; 
32'd10684: dataIn1 = 32'd10
; 
32'd10685: dataIn1 = 32'd11
; 
32'd10686: dataIn1 = 32'd12
; 
32'd10687: dataIn1 = 32'd14
; 
32'd10688: dataIn1 = 32'd15
; 
32'd10689: dataIn1 = 32'd16
; 
32'd10690: dataIn1 = 32'd17
; 
32'd10691: dataIn1 = 32'd18
; 
32'd10692: dataIn1 = 32'd19
; 
32'd10693: dataIn1 = 32'd21
; 
32'd10694: dataIn1 = 32'd23
; 
32'd10695: dataIn1 = 32'd24
; 
32'd10696: dataIn1 = 32'd25
; 
32'd10697: dataIn1 = 32'd26
; 
32'd10698: dataIn1 = 32'd27
; 
32'd10699: dataIn1 = 32'd28
; 
32'd10700: dataIn1 = 32'd29
; 
32'd10701: dataIn1 = 32'd30
; 
32'd10702: dataIn1 = 32'd31
; 
32'd10703: dataIn1 = 32'd; 
32'd10704: dataIn1 = 32'd; 
32'd10705: dataIn1 = 32'd; 
32'd10706: dataIn1 = 32'd; 
32'd10707: dataIn1 = 32'd; 
32'd10708: dataIn1 = 32'd; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd82; 
32'd3: dataIn2 = 32'd65; 
32'd4: dataIn2 = 32'd46; 
32'd5: dataIn2 = 32'd13; 
32'd6: dataIn2 = 32'd49; 
32'd7: dataIn2 = 32'd64; 
32'd8: dataIn2 = 32'd7; 
32'd9: dataIn2 = 32'd54; 
32'd10: dataIn2 = 32'd86; 
32'd11: dataIn2 = 32'd80; 
32'd12: dataIn2 = 32'd45; 
32'd13: dataIn2 = 32'd38; 
32'd14: dataIn2 = 32'd87; 
32'd15: dataIn2 = 32'd41; 
32'd16: dataIn2 = 32'd1; 
32'd17: dataIn2 = 32'd57; 
32'd18: dataIn2 = 32'd58; 
32'd19: dataIn2 = 32'd12; 
32'd20: dataIn2 = 32'd66; 
32'd21: dataIn2 = 32'd20; 
32'd22: dataIn2 = 32'd0; 
32'd23: dataIn2 = 32'd9; 
32'd24: dataIn2 = 32'd60; 
32'd25: dataIn2 = 32'd16; 
32'd26: dataIn2 = 32'd26; 
32'd27: dataIn2 = 32'd63; 
32'd28: dataIn2 = 32'd46; 
32'd29: dataIn2 = 32'd9; 
32'd30: dataIn2 = 32'd68; 
32'd31: dataIn2 = 32'd2; 
32'd32: dataIn2 = 32'd60; 
32'd33: dataIn2 = 32'd64; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd170: dataIn2 = 32'd3; 
32'd171: dataIn2 = 32'd23; 
32'd172: dataIn2 = 32'd13; 
32'd173: dataIn2 = 32'd51; 
32'd174: dataIn2 = 32'd23; 
32'd175: dataIn2 = 32'd36; 
32'd176: dataIn2 = 32'd64; 
32'd177: dataIn2 = 32'd44; 
32'd178: dataIn2 = 32'd9; 
32'd179: dataIn2 = 32'd33; 
32'd180: dataIn2 = 32'd56; 
32'd181: dataIn2 = 32'd42; 
32'd182: dataIn2 = 32'd65; 
32'd183: dataIn2 = 32'd83; 
32'd184: dataIn2 = 32'd22; 
32'd185: dataIn2 = 32'd74; 
32'd186: dataIn2 = 32'd53; 
32'd187: dataIn2 = 32'd17; 
32'd188: dataIn2 = 32'd30; 
32'd189: dataIn2 = 32'd69; 
32'd190: dataIn2 = 32'd84; 
32'd191: dataIn2 = 32'd19; 
32'd192: dataIn2 = 32'd80; 
32'd193: dataIn2 = 32'd26; 
32'd194: dataIn2 = 32'd71; 
32'd195: dataIn2 = 32'd18; 
32'd196: dataIn2 = 32'd75; 
32'd197: dataIn2 = 32'd91; 
32'd198: dataIn2 = 32'd48; 
32'd199: dataIn2 = 32'd35; 
32'd200: dataIn2 = 32'd99; 
32'd201: dataIn2 = 32'd77; 
32'd202: dataIn2 = 32'd53; 
32'd203: dataIn2 = 32'd17; 
32'd204: dataIn2 = 32'd94; 
32'd205: dataIn2 = 32'd72; 
32'd206: dataIn2 = 32'd19; 
32'd207: dataIn2 = 32'd4; 
32'd208: dataIn2 = 32'd29; 
32'd209: dataIn2 = 32'd40; 
32'd210: dataIn2 = 32'd80; 
32'd211: dataIn2 = 32'd59; 
32'd212: dataIn2 = 32'd58; 
32'd213: dataIn2 = 32'd93; 
32'd214: dataIn2 = 32'd7; 
32'd215: dataIn2 = 32'd97; 
32'd216: dataIn2 = 32'd82; 
32'd217: dataIn2 = 32'd44; 
32'd218: dataIn2 = 32'd65; 
32'd219: dataIn2 = 32'd43; 
32'd220: dataIn2 = 32'd92; 
32'd221: dataIn2 = 32'd24; 
32'd222: dataIn2 = 32'd43; 
32'd223: dataIn2 = 32'd64; 
32'd224: dataIn2 = 32'd64; 
32'd225: dataIn2 = 32'd7; 
32'd226: dataIn2 = 32'd38; 
32'd227: dataIn2 = 32'd96; 
32'd228: dataIn2 = 32'd88; 
32'd229: dataIn2 = 32'd65; 
32'd230: dataIn2 = 32'd88; 
32'd231: dataIn2 = 32'd42; 
32'd232: dataIn2 = 32'd16; 
32'd233: dataIn2 = 32'd92; 
32'd234: dataIn2 = 32'd30; 
32'd235: dataIn2 = 32'd23; 
32'd236: dataIn2 = 32'd85; 
32'd237: dataIn2 = 32'd10; 
32'd238: dataIn2 = 32'd70; 
32'd239: dataIn2 = 32'd31; 
32'd240: dataIn2 = 32'd21; 
32'd241: dataIn2 = 32'd57; 
32'd242: dataIn2 = 32'd88; 
32'd243: dataIn2 = 32'd80; 
32'd244: dataIn2 = 32'd73; 
32'd245: dataIn2 = 32'd17; 
32'd246: dataIn2 = 32'd70; 
32'd247: dataIn2 = 32'd31; 
32'd248: dataIn2 = 32'd43; 
32'd249: dataIn2 = 32'd27; 
32'd250: dataIn2 = 32'd66; 
32'd251: dataIn2 = 32'd77; 
32'd252: dataIn2 = 32'd67; 
32'd253: dataIn2 = 32'd59; 
32'd254: dataIn2 = 32'd27; 
32'd255: dataIn2 = 32'd99; 
32'd256: dataIn2 = 32'd58; 
32'd257: dataIn2 = 32'd59; 
32'd258: dataIn2 = 32'd82; 
32'd259: dataIn2 = 32'd30; 
32'd260: dataIn2 = 32'd88; 
32'd261: dataIn2 = 32'd99; 
32'd262: dataIn2 = 32'd27; 
32'd263: dataIn2 = 32'd1; 
32'd264: dataIn2 = 32'd40; 
32'd265: dataIn2 = 32'd63; 
32'd266: dataIn2 = 32'd33; 
32'd267: dataIn2 = 32'd83; 
32'd268: dataIn2 = 32'd62; 
32'd269: dataIn2 = 32'd19; 
32'd270: dataIn2 = 32'd43; 
32'd271: dataIn2 = 32'd6; 
32'd272: dataIn2 = 32'd40; 
32'd273: dataIn2 = 32'd41; 
32'd274: dataIn2 = 32'd34; 
32'd275: dataIn2 = 32'd23; 
32'd276: dataIn2 = 32'd41; 
32'd277: dataIn2 = 32'd80; 
32'd278: dataIn2 = 32'd2; 
32'd279: dataIn2 = 32'd52; 
32'd280: dataIn2 = 32'd66; 
32'd281: dataIn2 = 32'd94; 
32'd282: dataIn2 = 32'd54; 
32'd283: dataIn2 = 32'd3; 
32'd284: dataIn2 = 32'd90; 
32'd285: dataIn2 = 32'd45; 
32'd286: dataIn2 = 32'd77; 
32'd287: dataIn2 = 32'd6; 
32'd288: dataIn2 = 32'd92; 
32'd289: dataIn2 = 32'd42; 
32'd290: dataIn2 = 32'd18; 
32'd291: dataIn2 = 32'd74; 
32'd292: dataIn2 = 32'd30; 
32'd293: dataIn2 = 32'd70; 
32'd294: dataIn2 = 32'd44; 
32'd295: dataIn2 = 32'd9; 
32'd296: dataIn2 = 32'd16; 
32'd297: dataIn2 = 32'd52; 
32'd298: dataIn2 = 32'd13; 
32'd299: dataIn2 = 32'd59; 
32'd300: dataIn2 = 32'd67; 
32'd301: dataIn2 = 32'd29; 
32'd302: dataIn2 = 32'd94; 
32'd303: dataIn2 = 32'd60; 
32'd304: dataIn2 = 32'd46; 
32'd305: dataIn2 = 32'd33; 
32'd306: dataIn2 = 32'd77; 
32'd307: dataIn2 = 32'd47; 
32'd308: dataIn2 = 32'd96; 
32'd309: dataIn2 = 32'd1; 
32'd310: dataIn2 = 32'd24; 
32'd311: dataIn2 = 32'd62; 
32'd312: dataIn2 = 32'd19; 
32'd313: dataIn2 = 32'd79; 
32'd314: dataIn2 = 32'd85; 
32'd315: dataIn2 = 32'd71; 
32'd316: dataIn2 = 32'd48; 
32'd317: dataIn2 = 32'd94; 
32'd318: dataIn2 = 32'd92; 
32'd319: dataIn2 = 32'd35; 
32'd320: dataIn2 = 32'd16; 
32'd321: dataIn2 = 32'd86; 
32'd322: dataIn2 = 32'd75; 
32'd323: dataIn2 = 32'd62; 
32'd324: dataIn2 = 32'd95; 
32'd325: dataIn2 = 32'd40; 
32'd326: dataIn2 = 32'd61; 
32'd327: dataIn2 = 32'd79; 
32'd328: dataIn2 = 32'd37; 
32'd329: dataIn2 = 32'd56; 
32'd330: dataIn2 = 32'd74; 
32'd331: dataIn2 = 32'd63; 
32'd332: dataIn2 = 32'd18; 
32'd333: dataIn2 = 32'd36; 
32'd334: dataIn2 = 32'd34; 
32'd335: dataIn2 = 32'd30; 
32'd336: dataIn2 = 32'd56; 
32'd337: dataIn2 = 32'd80; 
32'd338: dataIn2 = 32'd84; 
32'd339: dataIn2 = 32'd35; 
32'd340: dataIn2 = 32'd25; 
32'd341: dataIn2 = 32'd10; 
32'd342: dataIn2 = 32'd21; 
32'd343: dataIn2 = 32'd98; 
32'd344: dataIn2 = 32'd40; 
32'd345: dataIn2 = 32'd88; 
32'd346: dataIn2 = 32'd24; 
32'd347: dataIn2 = 32'd93; 
32'd348: dataIn2 = 32'd84; 
32'd349: dataIn2 = 32'd41; 
32'd350: dataIn2 = 32'd76; 
32'd351: dataIn2 = 32'd15; 
32'd352: dataIn2 = 32'd99; 
32'd353: dataIn2 = 32'd63; 
32'd354: dataIn2 = 32'd33; 
32'd355: dataIn2 = 32'd31; 
32'd356: dataIn2 = 32'd0; 
32'd357: dataIn2 = 32'd63; 
32'd358: dataIn2 = 32'd6; 
32'd359: dataIn2 = 32'd10; 
32'd360: dataIn2 = 32'd99; 
32'd361: dataIn2 = 32'd62; 
32'd362: dataIn2 = 32'd65; 
32'd363: dataIn2 = 32'd57; 
32'd364: dataIn2 = 32'd100; 
32'd365: dataIn2 = 32'd49; 
32'd366: dataIn2 = 32'd3; 
32'd367: dataIn2 = 32'd27; 
32'd368: dataIn2 = 32'd16; 
32'd369: dataIn2 = 32'd79; 
32'd370: dataIn2 = 32'd84; 
32'd371: dataIn2 = 32'd69; 
32'd372: dataIn2 = 32'd29; 
32'd373: dataIn2 = 32'd54; 
32'd374: dataIn2 = 32'd95; 
32'd375: dataIn2 = 32'd30; 
32'd376: dataIn2 = 32'd42; 
32'd377: dataIn2 = 32'd1; 
32'd378: dataIn2 = 32'd27; 
32'd379: dataIn2 = 32'd4; 
32'd380: dataIn2 = 32'd13; 
32'd381: dataIn2 = 32'd84; 
32'd382: dataIn2 = 32'd66; 
32'd383: dataIn2 = 32'd34; 
32'd384: dataIn2 = 32'd76; 
32'd385: dataIn2 = 32'd72; 
32'd386: dataIn2 = 32'd6; 
32'd387: dataIn2 = 32'd4; 
32'd388: dataIn2 = 32'd38; 
32'd389: dataIn2 = 32'd38; 
32'd390: dataIn2 = 32'd20; 
32'd391: dataIn2 = 32'd29; 
32'd392: dataIn2 = 32'd25; 
32'd393: dataIn2 = 32'd19; 
32'd394: dataIn2 = 32'd22; 
32'd395: dataIn2 = 32'd96; 
32'd396: dataIn2 = 32'd74; 
32'd397: dataIn2 = 32'd32; 
32'd398: dataIn2 = 32'd89; 
32'd399: dataIn2 = 32'd5; 
32'd400: dataIn2 = 32'd12; 
32'd401: dataIn2 = 32'd87; 
32'd402: dataIn2 = 32'd85; 
32'd403: dataIn2 = 32'd67; 
32'd404: dataIn2 = 32'd39; 
32'd405: dataIn2 = 32'd0; 
32'd406: dataIn2 = 32'd90; 
32'd407: dataIn2 = 32'd77; 
32'd408: dataIn2 = 32'd57; 
32'd409: dataIn2 = 32'd50; 
32'd410: dataIn2 = 32'd90; 
32'd411: dataIn2 = 32'd2; 
32'd412: dataIn2 = 32'd36; 
32'd413: dataIn2 = 32'd26; 
32'd414: dataIn2 = 32'd96; 
32'd415: dataIn2 = 32'd77; 
32'd416: dataIn2 = 32'd20; 
32'd417: dataIn2 = 32'd15; 
32'd418: dataIn2 = 32'd54; 
32'd419: dataIn2 = 32'd94; 
32'd420: dataIn2 = 32'd22; 
32'd421: dataIn2 = 32'd22; 
32'd422: dataIn2 = 32'd6; 
32'd423: dataIn2 = 32'd96; 
32'd424: dataIn2 = 32'd83; 
32'd425: dataIn2 = 32'd58; 
32'd426: dataIn2 = 32'd35; 
32'd427: dataIn2 = 32'd71; 
32'd428: dataIn2 = 32'd79; 
32'd429: dataIn2 = 32'd73; 
32'd430: dataIn2 = 32'd3; 
32'd431: dataIn2 = 32'd8; 
32'd432: dataIn2 = 32'd71; 
32'd433: dataIn2 = 32'd13; 
32'd434: dataIn2 = 32'd52; 
32'd435: dataIn2 = 32'd42; 
32'd436: dataIn2 = 32'd71; 
32'd437: dataIn2 = 32'd35; 
32'd438: dataIn2 = 32'd8; 
32'd439: dataIn2 = 32'd44; 
32'd440: dataIn2 = 32'd19; 
32'd441: dataIn2 = 32'd77; 
32'd442: dataIn2 = 32'd73; 
32'd443: dataIn2 = 32'd32; 
32'd444: dataIn2 = 32'd45; 
32'd445: dataIn2 = 32'd79; 
32'd446: dataIn2 = 32'd32; 
32'd447: dataIn2 = 32'd97; 
32'd448: dataIn2 = 32'd47; 
32'd449: dataIn2 = 32'd44; 
32'd450: dataIn2 = 32'd48; 
32'd451: dataIn2 = 32'd11; 
32'd452: dataIn2 = 32'd99; 
32'd453: dataIn2 = 32'd14; 
32'd454: dataIn2 = 32'd27; 
32'd455: dataIn2 = 32'd6; 
32'd456: dataIn2 = 32'd12; 
32'd457: dataIn2 = 32'd89; 
32'd458: dataIn2 = 32'd87; 
32'd459: dataIn2 = 32'd7; 
32'd460: dataIn2 = 32'd0; 
32'd461: dataIn2 = 32'd21; 
32'd462: dataIn2 = 32'd29; 
32'd463: dataIn2 = 32'd33; 
32'd464: dataIn2 = 32'd66; 
32'd465: dataIn2 = 32'd80; 
32'd466: dataIn2 = 32'd20; 
32'd467: dataIn2 = 32'd91; 
32'd468: dataIn2 = 32'd30; 
32'd469: dataIn2 = 32'd56; 
32'd470: dataIn2 = 32'd59; 
32'd471: dataIn2 = 32'd45; 
32'd472: dataIn2 = 32'd13; 
32'd473: dataIn2 = 32'd52; 
32'd474: dataIn2 = 32'd43; 
32'd475: dataIn2 = 32'd59; 
32'd476: dataIn2 = 32'd42; 
32'd477: dataIn2 = 32'd17; 
32'd478: dataIn2 = 32'd76; 
32'd479: dataIn2 = 32'd51; 
32'd480: dataIn2 = 32'd46; 
32'd481: dataIn2 = 32'd46; 
32'd482: dataIn2 = 32'd0; 
32'd483: dataIn2 = 32'd50; 
32'd484: dataIn2 = 32'd72; 
32'd485: dataIn2 = 32'd0; 
32'd486: dataIn2 = 32'd69; 
32'd487: dataIn2 = 32'd14; 
32'd488: dataIn2 = 32'd56; 
32'd489: dataIn2 = 32'd21; 
32'd490: dataIn2 = 32'd88; 
32'd491: dataIn2 = 32'd24; 
32'd492: dataIn2 = 32'd11; 
32'd493: dataIn2 = 32'd2; 
32'd494: dataIn2 = 32'd58; 
32'd495: dataIn2 = 32'd4; 
32'd496: dataIn2 = 32'd28; 
32'd497: dataIn2 = 32'd13; 
32'd498: dataIn2 = 32'd45; 
32'd499: dataIn2 = 32'd88; 
32'd500: dataIn2 = 32'd6; 
32'd501: dataIn2 = 32'd99; 
32'd502: dataIn2 = 32'd41; 
32'd503: dataIn2 = 32'd16; 
32'd504: dataIn2 = 32'd75; 
32'd505: dataIn2 = 32'd87; 
32'd506: dataIn2 = 32'd100; 
32'd507: dataIn2 = 32'd40; 
32'd508: dataIn2 = 32'd1; 
32'd509: dataIn2 = 32'd90; 
32'd510: dataIn2 = 32'd51; 
32'd511: dataIn2 = 32'd3; 
32'd512: dataIn2 = 32'd55; 
32'd513: dataIn2 = 32'd36; 
32'd514: dataIn2 = 32'd99; 
32'd515: dataIn2 = 32'd96; 
32'd516: dataIn2 = 32'd93; 
32'd517: dataIn2 = 32'd61; 
32'd518: dataIn2 = 32'd82; 
32'd519: dataIn2 = 32'd99; 
32'd520: dataIn2 = 32'd74; 
32'd521: dataIn2 = 32'd70; 
32'd522: dataIn2 = 32'd74; 
32'd523: dataIn2 = 32'd75; 
32'd524: dataIn2 = 32'd60; 
32'd525: dataIn2 = 32'd47; 
32'd526: dataIn2 = 32'd24; 
32'd527: dataIn2 = 32'd72; 
32'd528: dataIn2 = 32'd87; 
32'd529: dataIn2 = 32'd62; 
32'd530: dataIn2 = 32'd78; 
32'd531: dataIn2 = 32'd24; 
32'd532: dataIn2 = 32'd82; 
32'd533: dataIn2 = 32'd0; 
32'd534: dataIn2 = 32'd97; 
32'd535: dataIn2 = 32'd43; 
32'd536: dataIn2 = 32'd96; 
32'd537: dataIn2 = 32'd23; 
32'd538: dataIn2 = 32'd35; 
32'd539: dataIn2 = 32'd9; 
32'd540: dataIn2 = 32'd82; 
32'd541: dataIn2 = 32'd58; 
32'd542: dataIn2 = 32'd10; 
32'd543: dataIn2 = 32'd39; 
32'd544: dataIn2 = 32'd77; 
32'd545: dataIn2 = 32'd19; 
32'd546: dataIn2 = 32'd31; 
32'd547: dataIn2 = 32'd61; 
32'd548: dataIn2 = 32'd85; 
32'd549: dataIn2 = 32'd22; 
32'd550: dataIn2 = 32'd3; 
32'd551: dataIn2 = 32'd50; 
32'd552: dataIn2 = 32'd51; 
32'd553: dataIn2 = 32'd42; 
32'd554: dataIn2 = 32'd37; 
32'd555: dataIn2 = 32'd12; 
32'd556: dataIn2 = 32'd51; 
32'd557: dataIn2 = 32'd31; 
32'd558: dataIn2 = 32'd97; 
32'd559: dataIn2 = 32'd39; 
32'd560: dataIn2 = 32'd100; 
32'd561: dataIn2 = 32'd51; 
32'd562: dataIn2 = 32'd37; 
32'd563: dataIn2 = 32'd6; 
32'd564: dataIn2 = 32'd35; 
32'd565: dataIn2 = 32'd13; 
32'd566: dataIn2 = 32'd3; 
32'd567: dataIn2 = 32'd88; 
32'd568: dataIn2 = 32'd2; 
32'd569: dataIn2 = 32'd74; 
32'd570: dataIn2 = 32'd12; 
32'd571: dataIn2 = 32'd31; 
32'd572: dataIn2 = 32'd66; 
32'd573: dataIn2 = 32'd95; 
32'd574: dataIn2 = 32'd4; 
32'd575: dataIn2 = 32'd39; 
32'd576: dataIn2 = 32'd22; 
32'd577: dataIn2 = 32'd7; 
32'd578: dataIn2 = 32'd34; 
32'd579: dataIn2 = 32'd95; 
32'd580: dataIn2 = 32'd4; 
32'd581: dataIn2 = 32'd34; 
32'd582: dataIn2 = 32'd23; 
32'd583: dataIn2 = 32'd48; 
32'd584: dataIn2 = 32'd23; 
32'd585: dataIn2 = 32'd34; 
32'd586: dataIn2 = 32'd53; 
32'd587: dataIn2 = 32'd93; 
32'd588: dataIn2 = 32'd87; 
32'd589: dataIn2 = 32'd33; 
32'd590: dataIn2 = 32'd68; 
32'd591: dataIn2 = 32'd37; 
32'd592: dataIn2 = 32'd5; 
32'd593: dataIn2 = 32'd71; 
32'd594: dataIn2 = 32'd24; 
32'd595: dataIn2 = 32'd24; 
32'd596: dataIn2 = 32'd47; 
32'd597: dataIn2 = 32'd46; 
32'd598: dataIn2 = 32'd42; 
32'd599: dataIn2 = 32'd47; 
32'd600: dataIn2 = 32'd98; 
32'd601: dataIn2 = 32'd15; 
32'd602: dataIn2 = 32'd7; 
32'd603: dataIn2 = 32'd30; 
32'd604: dataIn2 = 32'd35; 
32'd605: dataIn2 = 32'd7; 
32'd606: dataIn2 = 32'd89; 
32'd607: dataIn2 = 32'd19; 
32'd608: dataIn2 = 32'd98; 
32'd609: dataIn2 = 32'd99; 
32'd610: dataIn2 = 32'd25; 
32'd611: dataIn2 = 32'd89; 
32'd612: dataIn2 = 32'd89; 
32'd613: dataIn2 = 32'd32; 
32'd614: dataIn2 = 32'd40; 
32'd615: dataIn2 = 32'd42; 
32'd616: dataIn2 = 32'd50; 
32'd617: dataIn2 = 32'd94; 
32'd618: dataIn2 = 32'd40; 
32'd619: dataIn2 = 32'd22; 
32'd620: dataIn2 = 32'd16; 
32'd621: dataIn2 = 32'd67; 
32'd622: dataIn2 = 32'd73; 
32'd623: dataIn2 = 32'd39; 
32'd624: dataIn2 = 32'd15; 
32'd625: dataIn2 = 32'd92; 
32'd626: dataIn2 = 32'd42; 
32'd627: dataIn2 = 32'd48; 
32'd628: dataIn2 = 32'd37; 
32'd629: dataIn2 = 32'd63; 
32'd630: dataIn2 = 32'd68; 
32'd631: dataIn2 = 32'd34; 
32'd632: dataIn2 = 32'd52; 
32'd633: dataIn2 = 32'd24; 
32'd634: dataIn2 = 32'd55; 
32'd635: dataIn2 = 32'd64; 
32'd636: dataIn2 = 32'd70; 
32'd637: dataIn2 = 32'd30; 
32'd638: dataIn2 = 32'd75; 
32'd639: dataIn2 = 32'd36; 
32'd640: dataIn2 = 32'd49; 
32'd641: dataIn2 = 32'd5; 
32'd642: dataIn2 = 32'd25; 
32'd643: dataIn2 = 32'd35; 
32'd644: dataIn2 = 32'd67; 
32'd645: dataIn2 = 32'd53; 
32'd646: dataIn2 = 32'd55; 
32'd647: dataIn2 = 32'd100; 
32'd648: dataIn2 = 32'd70; 
32'd649: dataIn2 = 32'd94; 
32'd650: dataIn2 = 32'd55; 
32'd651: dataIn2 = 32'd72; 
32'd652: dataIn2 = 32'd52; 
32'd653: dataIn2 = 32'd57; 
32'd654: dataIn2 = 32'd29; 
32'd655: dataIn2 = 32'd60; 
32'd656: dataIn2 = 32'd75; 
32'd657: dataIn2 = 32'd11; 
32'd658: dataIn2 = 32'd36; 
32'd659: dataIn2 = 32'd15; 
32'd660: dataIn2 = 32'd40; 
32'd661: dataIn2 = 32'd18; 
32'd662: dataIn2 = 32'd15; 
32'd663: dataIn2 = 32'd73; 
32'd664: dataIn2 = 32'd56; 
32'd665: dataIn2 = 32'd97; 
32'd666: dataIn2 = 32'd26; 
32'd667: dataIn2 = 32'd10; 
32'd668: dataIn2 = 32'd87; 
32'd669: dataIn2 = 32'd20; 
32'd670: dataIn2 = 32'd42; 
32'd671: dataIn2 = 32'd38; 
32'd672: dataIn2 = 32'd74; 
32'd673: dataIn2 = 32'd40; 
32'd674: dataIn2 = 32'd48; 
32'd675: dataIn2 = 32'd100; 
32'd676: dataIn2 = 32'd49; 
32'd677: dataIn2 = 32'd81; 
32'd678: dataIn2 = 32'd30; 
32'd679: dataIn2 = 32'd1; 
32'd680: dataIn2 = 32'd18; 
32'd681: dataIn2 = 32'd80; 
32'd682: dataIn2 = 32'd67; 
32'd683: dataIn2 = 32'd78; 
32'd684: dataIn2 = 32'd49; 
32'd685: dataIn2 = 32'd10; 
32'd686: dataIn2 = 32'd63; 
32'd687: dataIn2 = 32'd83; 
32'd688: dataIn2 = 32'd80; 
32'd689: dataIn2 = 32'd1; 
32'd690: dataIn2 = 32'd31; 
32'd691: dataIn2 = 32'd9; 
32'd692: dataIn2 = 32'd36; 
32'd693: dataIn2 = 32'd52; 
32'd694: dataIn2 = 32'd63; 
32'd695: dataIn2 = 32'd26; 
32'd696: dataIn2 = 32'd68; 
32'd697: dataIn2 = 32'd7; 
32'd698: dataIn2 = 32'd16; 
32'd699: dataIn2 = 32'd49; 
32'd700: dataIn2 = 32'd30; 
32'd701: dataIn2 = 32'd11; 
32'd702: dataIn2 = 32'd62; 
32'd703: dataIn2 = 32'd62; 
32'd704: dataIn2 = 32'd54; 
32'd705: dataIn2 = 32'd32; 
32'd706: dataIn2 = 32'd72; 
32'd707: dataIn2 = 32'd80; 
32'd708: dataIn2 = 32'd91; 
32'd709: dataIn2 = 32'd37; 
32'd710: dataIn2 = 32'd90; 
32'd711: dataIn2 = 32'd89; 
32'd712: dataIn2 = 32'd41; 
32'd713: dataIn2 = 32'd9; 
32'd714: dataIn2 = 32'd91; 
32'd715: dataIn2 = 32'd44; 
32'd716: dataIn2 = 32'd1; 
32'd717: dataIn2 = 32'd73; 
32'd718: dataIn2 = 32'd9; 
32'd719: dataIn2 = 32'd57; 
32'd720: dataIn2 = 32'd91; 
32'd721: dataIn2 = 32'd61; 
32'd722: dataIn2 = 32'd61; 
32'd723: dataIn2 = 32'd95; 
32'd724: dataIn2 = 32'd71; 
32'd725: dataIn2 = 32'd87; 
32'd726: dataIn2 = 32'd36; 
32'd727: dataIn2 = 32'd67; 
32'd728: dataIn2 = 32'd87; 
32'd729: dataIn2 = 32'd0; 
32'd730: dataIn2 = 32'd0; 
32'd731: dataIn2 = 32'd34; 
32'd732: dataIn2 = 32'd46; 
32'd733: dataIn2 = 32'd59; 
32'd734: dataIn2 = 32'd52; 
32'd735: dataIn2 = 32'd63; 
32'd736: dataIn2 = 32'd17; 
32'd737: dataIn2 = 32'd89; 
32'd738: dataIn2 = 32'd81; 
32'd739: dataIn2 = 32'd10; 
32'd740: dataIn2 = 32'd86; 
32'd741: dataIn2 = 32'd94; 
32'd742: dataIn2 = 32'd1; 
32'd743: dataIn2 = 32'd71; 
32'd744: dataIn2 = 32'd16; 
32'd745: dataIn2 = 32'd83; 
32'd746: dataIn2 = 32'd59; 
32'd747: dataIn2 = 32'd15; 
32'd748: dataIn2 = 32'd70; 
32'd749: dataIn2 = 32'd35; 
32'd750: dataIn2 = 32'd83; 
32'd751: dataIn2 = 32'd91; 
32'd752: dataIn2 = 32'd54; 
32'd753: dataIn2 = 32'd3; 
32'd754: dataIn2 = 32'd84; 
32'd755: dataIn2 = 32'd60; 
32'd756: dataIn2 = 32'd39; 
32'd757: dataIn2 = 32'd97; 
32'd758: dataIn2 = 32'd75; 
32'd759: dataIn2 = 32'd69; 
32'd760: dataIn2 = 32'd58; 
32'd761: dataIn2 = 32'd78; 
32'd762: dataIn2 = 32'd20; 
32'd763: dataIn2 = 32'd17; 
32'd764: dataIn2 = 32'd54; 
32'd765: dataIn2 = 32'd56; 
32'd766: dataIn2 = 32'd20; 
32'd767: dataIn2 = 32'd97; 
32'd768: dataIn2 = 32'd42; 
32'd769: dataIn2 = 32'd69; 
32'd770: dataIn2 = 32'd72; 
32'd771: dataIn2 = 32'd70; 
32'd772: dataIn2 = 32'd61; 
32'd773: dataIn2 = 32'd61; 
32'd774: dataIn2 = 32'd82; 
32'd775: dataIn2 = 32'd44; 
32'd776: dataIn2 = 32'd87; 
32'd777: dataIn2 = 32'd41; 
32'd778: dataIn2 = 32'd18; 
32'd779: dataIn2 = 32'd78; 
32'd780: dataIn2 = 32'd54; 
32'd781: dataIn2 = 32'd16; 
32'd782: dataIn2 = 32'd10; 
32'd783: dataIn2 = 32'd95; 
32'd784: dataIn2 = 32'd97; 
32'd785: dataIn2 = 32'd12; 
32'd786: dataIn2 = 32'd19; 
32'd787: dataIn2 = 32'd28; 
32'd788: dataIn2 = 32'd71; 
32'd789: dataIn2 = 32'd49; 
32'd790: dataIn2 = 32'd11; 
32'd791: dataIn2 = 32'd80; 
32'd792: dataIn2 = 32'd39; 
32'd793: dataIn2 = 32'd42; 
32'd794: dataIn2 = 32'd96; 
32'd795: dataIn2 = 32'd25; 
32'd796: dataIn2 = 32'd40; 
32'd797: dataIn2 = 32'd2; 
32'd798: dataIn2 = 32'd55; 
32'd799: dataIn2 = 32'd50; 
32'd800: dataIn2 = 32'd26; 
32'd801: dataIn2 = 32'd94; 
32'd802: dataIn2 = 32'd51; 
32'd803: dataIn2 = 32'd27; 
32'd804: dataIn2 = 32'd77; 
32'd805: dataIn2 = 32'd15; 
32'd806: dataIn2 = 32'd92; 
32'd807: dataIn2 = 32'd4; 
32'd808: dataIn2 = 32'd22; 
32'd809: dataIn2 = 32'd12; 
32'd810: dataIn2 = 32'd25; 
32'd811: dataIn2 = 32'd85; 
32'd812: dataIn2 = 32'd46; 
32'd813: dataIn2 = 32'd9; 
32'd814: dataIn2 = 32'd78; 
32'd815: dataIn2 = 32'd84; 
32'd816: dataIn2 = 32'd11; 
32'd817: dataIn2 = 32'd70; 
32'd818: dataIn2 = 32'd90; 
32'd819: dataIn2 = 32'd38; 
32'd820: dataIn2 = 32'd16; 
32'd821: dataIn2 = 32'd96; 
32'd822: dataIn2 = 32'd62; 
32'd823: dataIn2 = 32'd44; 
32'd824: dataIn2 = 32'd0; 
32'd825: dataIn2 = 32'd42; 
32'd826: dataIn2 = 32'd79; 
32'd827: dataIn2 = 32'd14; 
32'd828: dataIn2 = 32'd83; 
32'd829: dataIn2 = 32'd22; 
32'd830: dataIn2 = 32'd95; 
32'd831: dataIn2 = 32'd62; 
32'd832: dataIn2 = 32'd76; 
32'd833: dataIn2 = 32'd83; 
32'd834: dataIn2 = 32'd87; 
32'd835: dataIn2 = 32'd1; 
32'd836: dataIn2 = 32'd99; 
32'd837: dataIn2 = 32'd34; 
32'd838: dataIn2 = 32'd15; 
32'd839: dataIn2 = 32'd80; 
32'd840: dataIn2 = 32'd81; 
32'd841: dataIn2 = 32'd5; 
32'd842: dataIn2 = 32'd98; 
32'd843: dataIn2 = 32'd78; 
32'd844: dataIn2 = 32'd45; 
32'd845: dataIn2 = 32'd99; 
32'd846: dataIn2 = 32'd62; 
32'd847: dataIn2 = 32'd73; 
32'd848: dataIn2 = 32'd97; 
32'd849: dataIn2 = 32'd37; 
32'd850: dataIn2 = 32'd58; 
32'd851: dataIn2 = 32'd98; 
32'd852: dataIn2 = 32'd73; 
32'd853: dataIn2 = 32'd14; 
32'd854: dataIn2 = 32'd23; 
32'd855: dataIn2 = 32'd43; 
32'd856: dataIn2 = 32'd93; 
32'd857: dataIn2 = 32'd50; 
32'd858: dataIn2 = 32'd24; 
32'd859: dataIn2 = 32'd28; 
32'd860: dataIn2 = 32'd16; 
32'd861: dataIn2 = 32'd44; 
32'd862: dataIn2 = 32'd1; 
32'd863: dataIn2 = 32'd94; 
32'd864: dataIn2 = 32'd37; 
32'd865: dataIn2 = 32'd56; 
32'd866: dataIn2 = 32'd61; 
32'd867: dataIn2 = 32'd59; 
32'd868: dataIn2 = 32'd82; 
32'd869: dataIn2 = 32'd88; 
32'd870: dataIn2 = 32'd1; 
32'd871: dataIn2 = 32'd30; 
32'd872: dataIn2 = 32'd5; 
32'd873: dataIn2 = 32'd93; 
32'd874: dataIn2 = 32'd51; 
32'd875: dataIn2 = 32'd56; 
32'd876: dataIn2 = 32'd33; 
32'd877: dataIn2 = 32'd26; 
32'd878: dataIn2 = 32'd44; 
32'd879: dataIn2 = 32'd77; 
32'd880: dataIn2 = 32'd74; 
32'd881: dataIn2 = 32'd50; 
32'd882: dataIn2 = 32'd31; 
32'd883: dataIn2 = 32'd53; 
32'd884: dataIn2 = 32'd68; 
32'd885: dataIn2 = 32'd93; 
32'd886: dataIn2 = 32'd45; 
32'd887: dataIn2 = 32'd1; 
32'd888: dataIn2 = 32'd4; 
32'd889: dataIn2 = 32'd77; 
32'd890: dataIn2 = 32'd15; 
32'd891: dataIn2 = 32'd28; 
32'd892: dataIn2 = 32'd71; 
32'd893: dataIn2 = 32'd69; 
32'd894: dataIn2 = 32'd93; 
32'd895: dataIn2 = 32'd29; 
32'd896: dataIn2 = 32'd89; 
32'd897: dataIn2 = 32'd42; 
32'd898: dataIn2 = 32'd33; 
32'd899: dataIn2 = 32'd97; 
32'd900: dataIn2 = 32'd69; 
32'd901: dataIn2 = 32'd32; 
32'd902: dataIn2 = 32'd42; 
32'd903: dataIn2 = 32'd1; 
32'd904: dataIn2 = 32'd24; 
32'd905: dataIn2 = 32'd89; 
32'd906: dataIn2 = 32'd11; 
32'd907: dataIn2 = 32'd4; 
32'd908: dataIn2 = 32'd79; 
32'd909: dataIn2 = 32'd50; 
32'd910: dataIn2 = 32'd52; 
32'd911: dataIn2 = 32'd48; 
32'd912: dataIn2 = 32'd92; 
32'd913: dataIn2 = 32'd100; 
32'd914: dataIn2 = 32'd40; 
32'd915: dataIn2 = 32'd62; 
32'd916: dataIn2 = 32'd92; 
32'd917: dataIn2 = 32'd94; 
32'd918: dataIn2 = 32'd17; 
32'd919: dataIn2 = 32'd81; 
32'd920: dataIn2 = 32'd31; 
32'd921: dataIn2 = 32'd65; 
32'd922: dataIn2 = 32'd0; 
32'd923: dataIn2 = 32'd26; 
32'd924: dataIn2 = 32'd62; 
32'd925: dataIn2 = 32'd31; 
32'd926: dataIn2 = 32'd60; 
32'd927: dataIn2 = 32'd27; 
32'd928: dataIn2 = 32'd34; 
32'd929: dataIn2 = 32'd55; 
32'd930: dataIn2 = 32'd70; 
32'd931: dataIn2 = 32'd65; 
32'd932: dataIn2 = 32'd43; 
32'd933: dataIn2 = 32'd37; 
32'd934: dataIn2 = 32'd50; 
32'd935: dataIn2 = 32'd73; 
32'd936: dataIn2 = 32'd10; 
32'd937: dataIn2 = 32'd82; 
32'd938: dataIn2 = 32'd100; 
32'd939: dataIn2 = 32'd39; 
32'd940: dataIn2 = 32'd97; 
32'd941: dataIn2 = 32'd88; 
32'd942: dataIn2 = 32'd32; 
32'd943: dataIn2 = 32'd37; 
32'd944: dataIn2 = 32'd39; 
32'd945: dataIn2 = 32'd63; 
32'd946: dataIn2 = 32'd43; 
32'd947: dataIn2 = 32'd58; 
32'd948: dataIn2 = 32'd32; 
32'd949: dataIn2 = 32'd28; 
32'd950: dataIn2 = 32'd88; 
32'd951: dataIn2 = 32'd56; 
32'd952: dataIn2 = 32'd59; 
32'd953: dataIn2 = 32'd93; 
32'd954: dataIn2 = 32'd85; 
32'd955: dataIn2 = 32'd40; 
32'd956: dataIn2 = 32'd11; 
32'd957: dataIn2 = 32'd59; 
32'd958: dataIn2 = 32'd47; 
32'd959: dataIn2 = 32'd9; 
32'd960: dataIn2 = 32'd95; 
32'd961: dataIn2 = 32'd36; 
32'd962: dataIn2 = 32'd94; 
32'd963: dataIn2 = 32'd34; 
32'd964: dataIn2 = 32'd73; 
32'd965: dataIn2 = 32'd12; 
32'd966: dataIn2 = 32'd72; 
32'd967: dataIn2 = 32'd14; 
32'd968: dataIn2 = 32'd0; 
32'd969: dataIn2 = 32'd17; 
32'd970: dataIn2 = 32'd42; 
32'd971: dataIn2 = 32'd8; 
32'd972: dataIn2 = 32'd71; 
32'd973: dataIn2 = 32'd62; 
32'd974: dataIn2 = 32'd12; 
32'd975: dataIn2 = 32'd86; 
32'd976: dataIn2 = 32'd48; 
32'd977: dataIn2 = 32'd71; 
32'd978: dataIn2 = 32'd6; 
32'd979: dataIn2 = 32'd62; 
32'd980: dataIn2 = 32'd51; 
32'd981: dataIn2 = 32'd52; 
32'd982: dataIn2 = 32'd62; 
32'd983: dataIn2 = 32'd64; 
32'd984: dataIn2 = 32'd65; 
32'd985: dataIn2 = 32'd80; 
32'd986: dataIn2 = 32'd40; 
32'd987: dataIn2 = 32'd64; 
32'd988: dataIn2 = 32'd43; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_32_20.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
