//64x64 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 2458 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd330 ; 
  wdata_col_base = 32'd27880 ; 
  row_base = 32'd303380 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #261000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd303380: dataIn1 = 32'd0
; 
32'd303381: dataIn1 = 32'd28
; 
32'd303382: dataIn1 = 32'd59
; 
32'd303383: dataIn1 = 32'd97
; 
32'd303384: dataIn1 = 32'd132
; 
32'd303385: dataIn1 = 32'd168
; 
32'd303386: dataIn1 = 32'd205
; 
32'd303387: dataIn1 = 32'd245
; 
32'd303388: dataIn1 = 32'd283
; 
32'd303389: dataIn1 = 32'd314
; 
32'd303390: dataIn1 = 32'd351
; 
32'd303391: dataIn1 = 32'd379
; 
32'd303392: dataIn1 = 32'd416
; 
32'd303393: dataIn1 = 32'd449
; 
32'd303394: dataIn1 = 32'd486
; 
32'd303395: dataIn1 = 32'd525
; 
32'd303396: dataIn1 = 32'd564
; 
32'd303397: dataIn1 = 32'd594
; 
32'd303398: dataIn1 = 32'd630
; 
32'd303399: dataIn1 = 32'd668
; 
32'd303400: dataIn1 = 32'd705
; 
32'd303401: dataIn1 = 32'd745
; 
32'd303402: dataIn1 = 32'd780
; 
32'd303403: dataIn1 = 32'd810
; 
32'd303404: dataIn1 = 32'd844
; 
32'd303405: dataIn1 = 32'd878
; 
32'd303406: dataIn1 = 32'd912
; 
32'd303407: dataIn1 = 32'd942
; 
32'd303408: dataIn1 = 32'd983
; 
32'd303409: dataIn1 = 32'd1018
; 
32'd303410: dataIn1 = 32'd1062
; 
32'd303411: dataIn1 = 32'd1098
; 
32'd303412: dataIn1 = 32'd1130
; 
32'd303413: dataIn1 = 32'd1172
; 
32'd303414: dataIn1 = 32'd1209
; 
32'd303415: dataIn1 = 32'd1248
; 
32'd303416: dataIn1 = 32'd1282
; 
32'd303417: dataIn1 = 32'd1315
; 
32'd303418: dataIn1 = 32'd1359
; 
32'd303419: dataIn1 = 32'd1396
; 
32'd303420: dataIn1 = 32'd1427
; 
32'd303421: dataIn1 = 32'd1460
; 
32'd303422: dataIn1 = 32'd1498
; 
32'd303423: dataIn1 = 32'd1536
; 
32'd303424: dataIn1 = 32'd1568
; 
32'd303425: dataIn1 = 32'd1606
; 
32'd303426: dataIn1 = 32'd1646
; 
32'd303427: dataIn1 = 32'd1680
; 
32'd303428: dataIn1 = 32'd1710
; 
32'd303429: dataIn1 = 32'd1746
; 
32'd303430: dataIn1 = 32'd1783
; 
32'd303431: dataIn1 = 32'd1818
; 
32'd303432: dataIn1 = 32'd1851
; 
32'd303433: dataIn1 = 32'd1880
; 
32'd303434: dataIn1 = 32'd1914
; 
32'd303435: dataIn1 = 32'd1951
; 
32'd303436: dataIn1 = 32'd1993
; 
32'd303437: dataIn1 = 32'd2034
; 
32'd303438: dataIn1 = 32'd2071
; 
32'd303439: dataIn1 = 32'd2104
; 
32'd303440: dataIn1 = 32'd2141
; 
32'd303441: dataIn1 = 32'd2177
; 
32'd303442: dataIn1 = 32'd2214
; 
32'd303443: dataIn1 = 32'd2247
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd27880: dataIn1 = 32'd0
; 
32'd27881: dataIn1 = 32'd28
; 
32'd27882: dataIn1 = 32'd59
; 
32'd27883: dataIn1 = 32'd97
; 
32'd27884: dataIn1 = 32'd132
; 
32'd27885: dataIn1 = 32'd168
; 
32'd27886: dataIn1 = 32'd205
; 
32'd27887: dataIn1 = 32'd245
; 
32'd27888: dataIn1 = 32'd283
; 
32'd27889: dataIn1 = 32'd314
; 
32'd27890: dataIn1 = 32'd351
; 
32'd27891: dataIn1 = 32'd379
; 
32'd27892: dataIn1 = 32'd416
; 
32'd27893: dataIn1 = 32'd449
; 
32'd27894: dataIn1 = 32'd486
; 
32'd27895: dataIn1 = 32'd525
; 
32'd27896: dataIn1 = 32'd564
; 
32'd27897: dataIn1 = 32'd594
; 
32'd27898: dataIn1 = 32'd630
; 
32'd27899: dataIn1 = 32'd668
; 
32'd27900: dataIn1 = 32'd705
; 
32'd27901: dataIn1 = 32'd745
; 
32'd27902: dataIn1 = 32'd780
; 
32'd27903: dataIn1 = 32'd810
; 
32'd27904: dataIn1 = 32'd844
; 
32'd27905: dataIn1 = 32'd878
; 
32'd27906: dataIn1 = 32'd912
; 
32'd27907: dataIn1 = 32'd942
; 
32'd27908: dataIn1 = 32'd983
; 
32'd27909: dataIn1 = 32'd1018
; 
32'd27910: dataIn1 = 32'd1062
; 
32'd27911: dataIn1 = 32'd1098
; 
32'd27912: dataIn1 = 32'd1130
; 
32'd27913: dataIn1 = 32'd1172
; 
32'd27914: dataIn1 = 32'd1209
; 
32'd27915: dataIn1 = 32'd1248
; 
32'd27916: dataIn1 = 32'd1282
; 
32'd27917: dataIn1 = 32'd1315
; 
32'd27918: dataIn1 = 32'd1359
; 
32'd27919: dataIn1 = 32'd1396
; 
32'd27920: dataIn1 = 32'd1427
; 
32'd27921: dataIn1 = 32'd1460
; 
32'd27922: dataIn1 = 32'd1498
; 
32'd27923: dataIn1 = 32'd1536
; 
32'd27924: dataIn1 = 32'd1568
; 
32'd27925: dataIn1 = 32'd1606
; 
32'd27926: dataIn1 = 32'd1646
; 
32'd27927: dataIn1 = 32'd1680
; 
32'd27928: dataIn1 = 32'd1710
; 
32'd27929: dataIn1 = 32'd1746
; 
32'd27930: dataIn1 = 32'd1783
; 
32'd27931: dataIn1 = 32'd1818
; 
32'd27932: dataIn1 = 32'd1851
; 
32'd27933: dataIn1 = 32'd1880
; 
32'd27934: dataIn1 = 32'd1914
; 
32'd27935: dataIn1 = 32'd1951
; 
32'd27936: dataIn1 = 32'd1993
; 
32'd27937: dataIn1 = 32'd2034
; 
32'd27938: dataIn1 = 32'd2071
; 
32'd27939: dataIn1 = 32'd2104
; 
32'd27940: dataIn1 = 32'd2141
; 
32'd27941: dataIn1 = 32'd2177
; 
32'd27942: dataIn1 = 32'd2214
; 
32'd27943: dataIn1 = 32'd2247
; 
32'd27944: dataIn1 = 32'd2283
; 
32'd27945: dataIn1 = 32'd1
; 
32'd27946: dataIn1 = 32'd3
; 
32'd27947: dataIn1 = 32'd6
; 
32'd27948: dataIn1 = 32'd9
; 
32'd27949: dataIn1 = 32'd10
; 
32'd27950: dataIn1 = 32'd11
; 
32'd27951: dataIn1 = 32'd13
; 
32'd27952: dataIn1 = 32'd17
; 
32'd27953: dataIn1 = 32'd18
; 
32'd27954: dataIn1 = 32'd19
; 
32'd27955: dataIn1 = 32'd22
; 
32'd27956: dataIn1 = 32'd24
; 
32'd27957: dataIn1 = 32'd26
; 
32'd27958: dataIn1 = 32'd29
; 
32'd27959: dataIn1 = 32'd30
; 
32'd27960: dataIn1 = 32'd31
; 
32'd27961: dataIn1 = 32'd33
; 
32'd27962: dataIn1 = 32'd37
; 
32'd27963: dataIn1 = 32'd40
; 
32'd27964: dataIn1 = 32'd42
; 
32'd27965: dataIn1 = 32'd45
; 
32'd27966: dataIn1 = 32'd48
; 
32'd27967: dataIn1 = 32'd50
; 
32'd27968: dataIn1 = 32'd53
; 
32'd27969: dataIn1 = 32'd58
; 
32'd27970: dataIn1 = 32'd59
; 
32'd27971: dataIn1 = 32'd60
; 
32'd27972: dataIn1 = 32'd61
; 
32'd27973: dataIn1 = 32'd5
; 
32'd27974: dataIn1 = 32'd9
; 
32'd27975: dataIn1 = 32'd10
; 
32'd27976: dataIn1 = 32'd11
; 
32'd27977: dataIn1 = 32'd13
; 
32'd27978: dataIn1 = 32'd14
; 
32'd27979: dataIn1 = 32'd16
; 
32'd27980: dataIn1 = 32'd21
; 
32'd27981: dataIn1 = 32'd23
; 
32'd27982: dataIn1 = 32'd25
; 
32'd27983: dataIn1 = 32'd26
; 
32'd27984: dataIn1 = 32'd29
; 
32'd27985: dataIn1 = 32'd30
; 
32'd27986: dataIn1 = 32'd31
; 
32'd27987: dataIn1 = 32'd34
; 
32'd27988: dataIn1 = 32'd37
; 
32'd27989: dataIn1 = 32'd38
; 
32'd27990: dataIn1 = 32'd39
; 
32'd27991: dataIn1 = 32'd44
; 
32'd27992: dataIn1 = 32'd45
; 
32'd27993: dataIn1 = 32'd47
; 
32'd27994: dataIn1 = 32'd48
; 
32'd27995: dataIn1 = 32'd49
; 
32'd27996: dataIn1 = 32'd50
; 
32'd27997: dataIn1 = 32'd51
; 
32'd27998: dataIn1 = 32'd52
; 
32'd27999: dataIn1 = 32'd57
; 
32'd28000: dataIn1 = 32'd58
; 
32'd28001: dataIn1 = 32'd60
; 
32'd28002: dataIn1 = 32'd62
; 
32'd28003: dataIn1 = 32'd63
; 
32'd28004: dataIn1 = 32'd0
; 
32'd28005: dataIn1 = 32'd3
; 
32'd28006: dataIn1 = 32'd4
; 
32'd28007: dataIn1 = 32'd5
; 
32'd28008: dataIn1 = 32'd6
; 
32'd28009: dataIn1 = 32'd7
; 
32'd28010: dataIn1 = 32'd8
; 
32'd28011: dataIn1 = 32'd9
; 
32'd28012: dataIn1 = 32'd12
; 
32'd28013: dataIn1 = 32'd13
; 
32'd28014: dataIn1 = 32'd15
; 
32'd28015: dataIn1 = 32'd16
; 
32'd28016: dataIn1 = 32'd17
; 
32'd28017: dataIn1 = 32'd19
; 
32'd28018: dataIn1 = 32'd22
; 
32'd28019: dataIn1 = 32'd25
; 
32'd28020: dataIn1 = 32'd26
; 
32'd28021: dataIn1 = 32'd27
; 
32'd28022: dataIn1 = 32'd28
; 
32'd28023: dataIn1 = 32'd30
; 
32'd28024: dataIn1 = 32'd31
; 
32'd28025: dataIn1 = 32'd34
; 
32'd28026: dataIn1 = 32'd35
; 
32'd28027: dataIn1 = 32'd36
; 
32'd28028: dataIn1 = 32'd38
; 
32'd28029: dataIn1 = 32'd40
; 
32'd28030: dataIn1 = 32'd41
; 
32'd28031: dataIn1 = 32'd42
; 
32'd28032: dataIn1 = 32'd44
; 
32'd28033: dataIn1 = 32'd45
; 
32'd28034: dataIn1 = 32'd47
; 
32'd28035: dataIn1 = 32'd48
; 
32'd28036: dataIn1 = 32'd50
; 
32'd28037: dataIn1 = 32'd52
; 
32'd28038: dataIn1 = 32'd56
; 
32'd28039: dataIn1 = 32'd58
; 
32'd28040: dataIn1 = 32'd59
; 
32'd28041: dataIn1 = 32'd62
; 
32'd28042: dataIn1 = 32'd0
; 
32'd28043: dataIn1 = 32'd1
; 
32'd28044: dataIn1 = 32'd3
; 
32'd28045: dataIn1 = 32'd4
; 
32'd28046: dataIn1 = 32'd9
; 
32'd28047: dataIn1 = 32'd10
; 
32'd28048: dataIn1 = 32'd11
; 
32'd28049: dataIn1 = 32'd12
; 
32'd28050: dataIn1 = 32'd13
; 
32'd28051: dataIn1 = 32'd17
; 
32'd28052: dataIn1 = 32'd18
; 
32'd28053: dataIn1 = 32'd20
; 
32'd28054: dataIn1 = 32'd22
; 
32'd28055: dataIn1 = 32'd25
; 
32'd28056: dataIn1 = 32'd27
; 
32'd28057: dataIn1 = 32'd32
; 
32'd28058: dataIn1 = 32'd33
; 
32'd28059: dataIn1 = 32'd34
; 
32'd28060: dataIn1 = 32'd36
; 
32'd28061: dataIn1 = 32'd42
; 
32'd28062: dataIn1 = 32'd43
; 
32'd28063: dataIn1 = 32'd45
; 
32'd28064: dataIn1 = 32'd46
; 
32'd28065: dataIn1 = 32'd48
; 
32'd28066: dataIn1 = 32'd50
; 
32'd28067: dataIn1 = 32'd52
; 
32'd28068: dataIn1 = 32'd54
; 
32'd28069: dataIn1 = 32'd55
; 
32'd28070: dataIn1 = 32'd56
; 
32'd28071: dataIn1 = 32'd57
; 
32'd28072: dataIn1 = 32'd58
; 
32'd28073: dataIn1 = 32'd59
; 
32'd28074: dataIn1 = 32'd60
; 
32'd28075: dataIn1 = 32'd61
; 
32'd28076: dataIn1 = 32'd62
; 
32'd28077: dataIn1 = 32'd0
; 
32'd28078: dataIn1 = 32'd1
; 
32'd28079: dataIn1 = 32'd3
; 
32'd28080: dataIn1 = 32'd4
; 
32'd28081: dataIn1 = 32'd5
; 
32'd28082: dataIn1 = 32'd6
; 
32'd28083: dataIn1 = 32'd9
; 
32'd28084: dataIn1 = 32'd10
; 
32'd28085: dataIn1 = 32'd11
; 
32'd28086: dataIn1 = 32'd12
; 
32'd28087: dataIn1 = 32'd14
; 
32'd28088: dataIn1 = 32'd15
; 
32'd28089: dataIn1 = 32'd16
; 
32'd28090: dataIn1 = 32'd17
; 
32'd28091: dataIn1 = 32'd21
; 
32'd28092: dataIn1 = 32'd23
; 
32'd28093: dataIn1 = 32'd24
; 
32'd28094: dataIn1 = 32'd28
; 
32'd28095: dataIn1 = 32'd30
; 
32'd28096: dataIn1 = 32'd31
; 
32'd28097: dataIn1 = 32'd32
; 
32'd28098: dataIn1 = 32'd33
; 
32'd28099: dataIn1 = 32'd34
; 
32'd28100: dataIn1 = 32'd36
; 
32'd28101: dataIn1 = 32'd41
; 
32'd28102: dataIn1 = 32'd42
; 
32'd28103: dataIn1 = 32'd43
; 
32'd28104: dataIn1 = 32'd44
; 
32'd28105: dataIn1 = 32'd46
; 
32'd28106: dataIn1 = 32'd47
; 
32'd28107: dataIn1 = 32'd48
; 
32'd28108: dataIn1 = 32'd49
; 
32'd28109: dataIn1 = 32'd50
; 
32'd28110: dataIn1 = 32'd52
; 
32'd28111: dataIn1 = 32'd54
; 
32'd28112: dataIn1 = 32'd61
; 
32'd28113: dataIn1 = 32'd0
; 
32'd28114: dataIn1 = 32'd2
; 
32'd28115: dataIn1 = 32'd3
; 
32'd28116: dataIn1 = 32'd5
; 
32'd28117: dataIn1 = 32'd6
; 
32'd28118: dataIn1 = 32'd7
; 
32'd28119: dataIn1 = 32'd8
; 
32'd28120: dataIn1 = 32'd9
; 
32'd28121: dataIn1 = 32'd10
; 
32'd28122: dataIn1 = 32'd11
; 
32'd28123: dataIn1 = 32'd13
; 
32'd28124: dataIn1 = 32'd17
; 
32'd28125: dataIn1 = 32'd18
; 
32'd28126: dataIn1 = 32'd19
; 
32'd28127: dataIn1 = 32'd21
; 
32'd28128: dataIn1 = 32'd22
; 
32'd28129: dataIn1 = 32'd24
; 
32'd28130: dataIn1 = 32'd25
; 
32'd28131: dataIn1 = 32'd26
; 
32'd28132: dataIn1 = 32'd27
; 
32'd28133: dataIn1 = 32'd28
; 
32'd28134: dataIn1 = 32'd30
; 
32'd28135: dataIn1 = 32'd34
; 
32'd28136: dataIn1 = 32'd36
; 
32'd28137: dataIn1 = 32'd39
; 
32'd28138: dataIn1 = 32'd41
; 
32'd28139: dataIn1 = 32'd42
; 
32'd28140: dataIn1 = 32'd43
; 
32'd28141: dataIn1 = 32'd44
; 
32'd28142: dataIn1 = 32'd45
; 
32'd28143: dataIn1 = 32'd46
; 
32'd28144: dataIn1 = 32'd50
; 
32'd28145: dataIn1 = 32'd55
; 
32'd28146: dataIn1 = 32'd58
; 
32'd28147: dataIn1 = 32'd60
; 
32'd28148: dataIn1 = 32'd61
; 
32'd28149: dataIn1 = 32'd63
; 
32'd28150: dataIn1 = 32'd0
; 
32'd28151: dataIn1 = 32'd1
; 
32'd28152: dataIn1 = 32'd2
; 
32'd28153: dataIn1 = 32'd3
; 
32'd28154: dataIn1 = 32'd9
; 
32'd28155: dataIn1 = 32'd10
; 
32'd28156: dataIn1 = 32'd11
; 
32'd28157: dataIn1 = 32'd12
; 
32'd28158: dataIn1 = 32'd13
; 
32'd28159: dataIn1 = 32'd14
; 
32'd28160: dataIn1 = 32'd15
; 
32'd28161: dataIn1 = 32'd17
; 
32'd28162: dataIn1 = 32'd18
; 
32'd28163: dataIn1 = 32'd19
; 
32'd28164: dataIn1 = 32'd21
; 
32'd28165: dataIn1 = 32'd22
; 
32'd28166: dataIn1 = 32'd26
; 
32'd28167: dataIn1 = 32'd27
; 
32'd28168: dataIn1 = 32'd28
; 
32'd28169: dataIn1 = 32'd29
; 
32'd28170: dataIn1 = 32'd30
; 
32'd28171: dataIn1 = 32'd31
; 
32'd28172: dataIn1 = 32'd32
; 
32'd28173: dataIn1 = 32'd33
; 
32'd28174: dataIn1 = 32'd36
; 
32'd28175: dataIn1 = 32'd37
; 
32'd28176: dataIn1 = 32'd38
; 
32'd28177: dataIn1 = 32'd40
; 
32'd28178: dataIn1 = 32'd42
; 
32'd28179: dataIn1 = 32'd43
; 
32'd28180: dataIn1 = 32'd46
; 
32'd28181: dataIn1 = 32'd47
; 
32'd28182: dataIn1 = 32'd50
; 
32'd28183: dataIn1 = 32'd52
; 
32'd28184: dataIn1 = 32'd55
; 
32'd28185: dataIn1 = 32'd56
; 
32'd28186: dataIn1 = 32'd57
; 
32'd28187: dataIn1 = 32'd59
; 
32'd28188: dataIn1 = 32'd60
; 
32'd28189: dataIn1 = 32'd63
; 
32'd28190: dataIn1 = 32'd3
; 
32'd28191: dataIn1 = 32'd6
; 
32'd28192: dataIn1 = 32'd8
; 
32'd28193: dataIn1 = 32'd9
; 
32'd28194: dataIn1 = 32'd11
; 
32'd28195: dataIn1 = 32'd12
; 
32'd28196: dataIn1 = 32'd14
; 
32'd28197: dataIn1 = 32'd15
; 
32'd28198: dataIn1 = 32'd16
; 
32'd28199: dataIn1 = 32'd17
; 
32'd28200: dataIn1 = 32'd19
; 
32'd28201: dataIn1 = 32'd20
; 
32'd28202: dataIn1 = 32'd22
; 
32'd28203: dataIn1 = 32'd24
; 
32'd28204: dataIn1 = 32'd26
; 
32'd28205: dataIn1 = 32'd27
; 
32'd28206: dataIn1 = 32'd28
; 
32'd28207: dataIn1 = 32'd31
; 
32'd28208: dataIn1 = 32'd32
; 
32'd28209: dataIn1 = 32'd33
; 
32'd28210: dataIn1 = 32'd35
; 
32'd28211: dataIn1 = 32'd37
; 
32'd28212: dataIn1 = 32'd38
; 
32'd28213: dataIn1 = 32'd39
; 
32'd28214: dataIn1 = 32'd40
; 
32'd28215: dataIn1 = 32'd41
; 
32'd28216: dataIn1 = 32'd44
; 
32'd28217: dataIn1 = 32'd45
; 
32'd28218: dataIn1 = 32'd46
; 
32'd28219: dataIn1 = 32'd47
; 
32'd28220: dataIn1 = 32'd48
; 
32'd28221: dataIn1 = 32'd49
; 
32'd28222: dataIn1 = 32'd50
; 
32'd28223: dataIn1 = 32'd51
; 
32'd28224: dataIn1 = 32'd52
; 
32'd28225: dataIn1 = 32'd54
; 
32'd28226: dataIn1 = 32'd57
; 
32'd28227: dataIn1 = 32'd58
; 
32'd28228: dataIn1 = 32'd3
; 
32'd28229: dataIn1 = 32'd4
; 
32'd28230: dataIn1 = 32'd5
; 
32'd28231: dataIn1 = 32'd6
; 
32'd28232: dataIn1 = 32'd7
; 
32'd28233: dataIn1 = 32'd9
; 
32'd28234: dataIn1 = 32'd11
; 
32'd28235: dataIn1 = 32'd13
; 
32'd28236: dataIn1 = 32'd19
; 
32'd28237: dataIn1 = 32'd25
; 
32'd28238: dataIn1 = 32'd26
; 
32'd28239: dataIn1 = 32'd27
; 
32'd28240: dataIn1 = 32'd28
; 
32'd28241: dataIn1 = 32'd32
; 
32'd28242: dataIn1 = 32'd33
; 
32'd28243: dataIn1 = 32'd36
; 
32'd28244: dataIn1 = 32'd37
; 
32'd28245: dataIn1 = 32'd38
; 
32'd28246: dataIn1 = 32'd40
; 
32'd28247: dataIn1 = 32'd41
; 
32'd28248: dataIn1 = 32'd42
; 
32'd28249: dataIn1 = 32'd45
; 
32'd28250: dataIn1 = 32'd47
; 
32'd28251: dataIn1 = 32'd48
; 
32'd28252: dataIn1 = 32'd49
; 
32'd28253: dataIn1 = 32'd50
; 
32'd28254: dataIn1 = 32'd51
; 
32'd28255: dataIn1 = 32'd53
; 
32'd28256: dataIn1 = 32'd54
; 
32'd28257: dataIn1 = 32'd60
; 
32'd28258: dataIn1 = 32'd63
; 
32'd28259: dataIn1 = 32'd0
; 
32'd28260: dataIn1 = 32'd1
; 
32'd28261: dataIn1 = 32'd2
; 
32'd28262: dataIn1 = 32'd4
; 
32'd28263: dataIn1 = 32'd7
; 
32'd28264: dataIn1 = 32'd8
; 
32'd28265: dataIn1 = 32'd9
; 
32'd28266: dataIn1 = 32'd10
; 
32'd28267: dataIn1 = 32'd11
; 
32'd28268: dataIn1 = 32'd13
; 
32'd28269: dataIn1 = 32'd14
; 
32'd28270: dataIn1 = 32'd15
; 
32'd28271: dataIn1 = 32'd17
; 
32'd28272: dataIn1 = 32'd20
; 
32'd28273: dataIn1 = 32'd21
; 
32'd28274: dataIn1 = 32'd23
; 
32'd28275: dataIn1 = 32'd24
; 
32'd28276: dataIn1 = 32'd26
; 
32'd28277: dataIn1 = 32'd28
; 
32'd28278: dataIn1 = 32'd34
; 
32'd28279: dataIn1 = 32'd36
; 
32'd28280: dataIn1 = 32'd37
; 
32'd28281: dataIn1 = 32'd39
; 
32'd28282: dataIn1 = 32'd40
; 
32'd28283: dataIn1 = 32'd41
; 
32'd28284: dataIn1 = 32'd42
; 
32'd28285: dataIn1 = 32'd43
; 
32'd28286: dataIn1 = 32'd44
; 
32'd28287: dataIn1 = 32'd51
; 
32'd28288: dataIn1 = 32'd52
; 
32'd28289: dataIn1 = 32'd53
; 
32'd28290: dataIn1 = 32'd56
; 
32'd28291: dataIn1 = 32'd57
; 
32'd28292: dataIn1 = 32'd58
; 
32'd28293: dataIn1 = 32'd59
; 
32'd28294: dataIn1 = 32'd61
; 
32'd28295: dataIn1 = 32'd62
; 
32'd28296: dataIn1 = 32'd1
; 
32'd28297: dataIn1 = 32'd2
; 
32'd28298: dataIn1 = 32'd5
; 
32'd28299: dataIn1 = 32'd8
; 
32'd28300: dataIn1 = 32'd10
; 
32'd28301: dataIn1 = 32'd18
; 
32'd28302: dataIn1 = 32'd19
; 
32'd28303: dataIn1 = 32'd23
; 
32'd28304: dataIn1 = 32'd25
; 
32'd28305: dataIn1 = 32'd27
; 
32'd28306: dataIn1 = 32'd28
; 
32'd28307: dataIn1 = 32'd31
; 
32'd28308: dataIn1 = 32'd33
; 
32'd28309: dataIn1 = 32'd35
; 
32'd28310: dataIn1 = 32'd36
; 
32'd28311: dataIn1 = 32'd37
; 
32'd28312: dataIn1 = 32'd40
; 
32'd28313: dataIn1 = 32'd44
; 
32'd28314: dataIn1 = 32'd46
; 
32'd28315: dataIn1 = 32'd47
; 
32'd28316: dataIn1 = 32'd48
; 
32'd28317: dataIn1 = 32'd50
; 
32'd28318: dataIn1 = 32'd51
; 
32'd28319: dataIn1 = 32'd55
; 
32'd28320: dataIn1 = 32'd56
; 
32'd28321: dataIn1 = 32'd58
; 
32'd28322: dataIn1 = 32'd60
; 
32'd28323: dataIn1 = 32'd61
; 
32'd28324: dataIn1 = 32'd1
; 
32'd28325: dataIn1 = 32'd2
; 
32'd28326: dataIn1 = 32'd3
; 
32'd28327: dataIn1 = 32'd4
; 
32'd28328: dataIn1 = 32'd8
; 
32'd28329: dataIn1 = 32'd10
; 
32'd28330: dataIn1 = 32'd11
; 
32'd28331: dataIn1 = 32'd12
; 
32'd28332: dataIn1 = 32'd13
; 
32'd28333: dataIn1 = 32'd14
; 
32'd28334: dataIn1 = 32'd15
; 
32'd28335: dataIn1 = 32'd16
; 
32'd28336: dataIn1 = 32'd17
; 
32'd28337: dataIn1 = 32'd19
; 
32'd28338: dataIn1 = 32'd23
; 
32'd28339: dataIn1 = 32'd25
; 
32'd28340: dataIn1 = 32'd26
; 
32'd28341: dataIn1 = 32'd29
; 
32'd28342: dataIn1 = 32'd31
; 
32'd28343: dataIn1 = 32'd32
; 
32'd28344: dataIn1 = 32'd36
; 
32'd28345: dataIn1 = 32'd37
; 
32'd28346: dataIn1 = 32'd39
; 
32'd28347: dataIn1 = 32'd40
; 
32'd28348: dataIn1 = 32'd42
; 
32'd28349: dataIn1 = 32'd43
; 
32'd28350: dataIn1 = 32'd44
; 
32'd28351: dataIn1 = 32'd46
; 
32'd28352: dataIn1 = 32'd47
; 
32'd28353: dataIn1 = 32'd51
; 
32'd28354: dataIn1 = 32'd53
; 
32'd28355: dataIn1 = 32'd54
; 
32'd28356: dataIn1 = 32'd57
; 
32'd28357: dataIn1 = 32'd58
; 
32'd28358: dataIn1 = 32'd61
; 
32'd28359: dataIn1 = 32'd62
; 
32'd28360: dataIn1 = 32'd63
; 
32'd28361: dataIn1 = 32'd1
; 
32'd28362: dataIn1 = 32'd2
; 
32'd28363: dataIn1 = 32'd4
; 
32'd28364: dataIn1 = 32'd5
; 
32'd28365: dataIn1 = 32'd6
; 
32'd28366: dataIn1 = 32'd7
; 
32'd28367: dataIn1 = 32'd13
; 
32'd28368: dataIn1 = 32'd14
; 
32'd28369: dataIn1 = 32'd16
; 
32'd28370: dataIn1 = 32'd20
; 
32'd28371: dataIn1 = 32'd23
; 
32'd28372: dataIn1 = 32'd24
; 
32'd28373: dataIn1 = 32'd27
; 
32'd28374: dataIn1 = 32'd28
; 
32'd28375: dataIn1 = 32'd31
; 
32'd28376: dataIn1 = 32'd32
; 
32'd28377: dataIn1 = 32'd33
; 
32'd28378: dataIn1 = 32'd34
; 
32'd28379: dataIn1 = 32'd35
; 
32'd28380: dataIn1 = 32'd37
; 
32'd28381: dataIn1 = 32'd39
; 
32'd28382: dataIn1 = 32'd41
; 
32'd28383: dataIn1 = 32'd43
; 
32'd28384: dataIn1 = 32'd44
; 
32'd28385: dataIn1 = 32'd46
; 
32'd28386: dataIn1 = 32'd51
; 
32'd28387: dataIn1 = 32'd52
; 
32'd28388: dataIn1 = 32'd56
; 
32'd28389: dataIn1 = 32'd57
; 
32'd28390: dataIn1 = 32'd59
; 
32'd28391: dataIn1 = 32'd61
; 
32'd28392: dataIn1 = 32'd62
; 
32'd28393: dataIn1 = 32'd63
; 
32'd28394: dataIn1 = 32'd0
; 
32'd28395: dataIn1 = 32'd4
; 
32'd28396: dataIn1 = 32'd5
; 
32'd28397: dataIn1 = 32'd9
; 
32'd28398: dataIn1 = 32'd10
; 
32'd28399: dataIn1 = 32'd12
; 
32'd28400: dataIn1 = 32'd13
; 
32'd28401: dataIn1 = 32'd15
; 
32'd28402: dataIn1 = 32'd16
; 
32'd28403: dataIn1 = 32'd17
; 
32'd28404: dataIn1 = 32'd18
; 
32'd28405: dataIn1 = 32'd20
; 
32'd28406: dataIn1 = 32'd25
; 
32'd28407: dataIn1 = 32'd27
; 
32'd28408: dataIn1 = 32'd28
; 
32'd28409: dataIn1 = 32'd29
; 
32'd28410: dataIn1 = 32'd30
; 
32'd28411: dataIn1 = 32'd31
; 
32'd28412: dataIn1 = 32'd33
; 
32'd28413: dataIn1 = 32'd35
; 
32'd28414: dataIn1 = 32'd37
; 
32'd28415: dataIn1 = 32'd38
; 
32'd28416: dataIn1 = 32'd41
; 
32'd28417: dataIn1 = 32'd42
; 
32'd28418: dataIn1 = 32'd43
; 
32'd28419: dataIn1 = 32'd44
; 
32'd28420: dataIn1 = 32'd45
; 
32'd28421: dataIn1 = 32'd46
; 
32'd28422: dataIn1 = 32'd51
; 
32'd28423: dataIn1 = 32'd53
; 
32'd28424: dataIn1 = 32'd55
; 
32'd28425: dataIn1 = 32'd56
; 
32'd28426: dataIn1 = 32'd58
; 
32'd28427: dataIn1 = 32'd59
; 
32'd28428: dataIn1 = 32'd60
; 
32'd28429: dataIn1 = 32'd61
; 
32'd28430: dataIn1 = 32'd62
; 
32'd28431: dataIn1 = 32'd0
; 
32'd28432: dataIn1 = 32'd1
; 
32'd28433: dataIn1 = 32'd2
; 
32'd28434: dataIn1 = 32'd3
; 
32'd28435: dataIn1 = 32'd4
; 
32'd28436: dataIn1 = 32'd5
; 
32'd28437: dataIn1 = 32'd7
; 
32'd28438: dataIn1 = 32'd8
; 
32'd28439: dataIn1 = 32'd13
; 
32'd28440: dataIn1 = 32'd15
; 
32'd28441: dataIn1 = 32'd16
; 
32'd28442: dataIn1 = 32'd18
; 
32'd28443: dataIn1 = 32'd20
; 
32'd28444: dataIn1 = 32'd22
; 
32'd28445: dataIn1 = 32'd25
; 
32'd28446: dataIn1 = 32'd26
; 
32'd28447: dataIn1 = 32'd28
; 
32'd28448: dataIn1 = 32'd30
; 
32'd28449: dataIn1 = 32'd31
; 
32'd28450: dataIn1 = 32'd32
; 
32'd28451: dataIn1 = 32'd33
; 
32'd28452: dataIn1 = 32'd36
; 
32'd28453: dataIn1 = 32'd37
; 
32'd28454: dataIn1 = 32'd38
; 
32'd28455: dataIn1 = 32'd40
; 
32'd28456: dataIn1 = 32'd41
; 
32'd28457: dataIn1 = 32'd43
; 
32'd28458: dataIn1 = 32'd46
; 
32'd28459: dataIn1 = 32'd47
; 
32'd28460: dataIn1 = 32'd48
; 
32'd28461: dataIn1 = 32'd49
; 
32'd28462: dataIn1 = 32'd50
; 
32'd28463: dataIn1 = 32'd51
; 
32'd28464: dataIn1 = 32'd54
; 
32'd28465: dataIn1 = 32'd55
; 
32'd28466: dataIn1 = 32'd56
; 
32'd28467: dataIn1 = 32'd57
; 
32'd28468: dataIn1 = 32'd60
; 
32'd28469: dataIn1 = 32'd61
; 
32'd28470: dataIn1 = 32'd0
; 
32'd28471: dataIn1 = 32'd1
; 
32'd28472: dataIn1 = 32'd7
; 
32'd28473: dataIn1 = 32'd8
; 
32'd28474: dataIn1 = 32'd9
; 
32'd28475: dataIn1 = 32'd11
; 
32'd28476: dataIn1 = 32'd12
; 
32'd28477: dataIn1 = 32'd14
; 
32'd28478: dataIn1 = 32'd15
; 
32'd28479: dataIn1 = 32'd16
; 
32'd28480: dataIn1 = 32'd18
; 
32'd28481: dataIn1 = 32'd19
; 
32'd28482: dataIn1 = 32'd20
; 
32'd28483: dataIn1 = 32'd21
; 
32'd28484: dataIn1 = 32'd22
; 
32'd28485: dataIn1 = 32'd23
; 
32'd28486: dataIn1 = 32'd25
; 
32'd28487: dataIn1 = 32'd27
; 
32'd28488: dataIn1 = 32'd28
; 
32'd28489: dataIn1 = 32'd29
; 
32'd28490: dataIn1 = 32'd30
; 
32'd28491: dataIn1 = 32'd32
; 
32'd28492: dataIn1 = 32'd33
; 
32'd28493: dataIn1 = 32'd35
; 
32'd28494: dataIn1 = 32'd36
; 
32'd28495: dataIn1 = 32'd38
; 
32'd28496: dataIn1 = 32'd41
; 
32'd28497: dataIn1 = 32'd42
; 
32'd28498: dataIn1 = 32'd44
; 
32'd28499: dataIn1 = 32'd47
; 
32'd28500: dataIn1 = 32'd48
; 
32'd28501: dataIn1 = 32'd49
; 
32'd28502: dataIn1 = 32'd51
; 
32'd28503: dataIn1 = 32'd53
; 
32'd28504: dataIn1 = 32'd54
; 
32'd28505: dataIn1 = 32'd57
; 
32'd28506: dataIn1 = 32'd59
; 
32'd28507: dataIn1 = 32'd60
; 
32'd28508: dataIn1 = 32'd63
; 
32'd28509: dataIn1 = 32'd0
; 
32'd28510: dataIn1 = 32'd3
; 
32'd28511: dataIn1 = 32'd7
; 
32'd28512: dataIn1 = 32'd9
; 
32'd28513: dataIn1 = 32'd10
; 
32'd28514: dataIn1 = 32'd11
; 
32'd28515: dataIn1 = 32'd14
; 
32'd28516: dataIn1 = 32'd15
; 
32'd28517: dataIn1 = 32'd16
; 
32'd28518: dataIn1 = 32'd20
; 
32'd28519: dataIn1 = 32'd22
; 
32'd28520: dataIn1 = 32'd24
; 
32'd28521: dataIn1 = 32'd25
; 
32'd28522: dataIn1 = 32'd26
; 
32'd28523: dataIn1 = 32'd28
; 
32'd28524: dataIn1 = 32'd31
; 
32'd28525: dataIn1 = 32'd32
; 
32'd28526: dataIn1 = 32'd36
; 
32'd28527: dataIn1 = 32'd37
; 
32'd28528: dataIn1 = 32'd38
; 
32'd28529: dataIn1 = 32'd40
; 
32'd28530: dataIn1 = 32'd41
; 
32'd28531: dataIn1 = 32'd43
; 
32'd28532: dataIn1 = 32'd47
; 
32'd28533: dataIn1 = 32'd51
; 
32'd28534: dataIn1 = 32'd53
; 
32'd28535: dataIn1 = 32'd55
; 
32'd28536: dataIn1 = 32'd56
; 
32'd28537: dataIn1 = 32'd57
; 
32'd28538: dataIn1 = 32'd61
; 
32'd28539: dataIn1 = 32'd1
; 
32'd28540: dataIn1 = 32'd4
; 
32'd28541: dataIn1 = 32'd6
; 
32'd28542: dataIn1 = 32'd10
; 
32'd28543: dataIn1 = 32'd12
; 
32'd28544: dataIn1 = 32'd13
; 
32'd28545: dataIn1 = 32'd16
; 
32'd28546: dataIn1 = 32'd22
; 
32'd28547: dataIn1 = 32'd24
; 
32'd28548: dataIn1 = 32'd25
; 
32'd28549: dataIn1 = 32'd26
; 
32'd28550: dataIn1 = 32'd28
; 
32'd28551: dataIn1 = 32'd29
; 
32'd28552: dataIn1 = 32'd30
; 
32'd28553: dataIn1 = 32'd31
; 
32'd28554: dataIn1 = 32'd32
; 
32'd28555: dataIn1 = 32'd33
; 
32'd28556: dataIn1 = 32'd34
; 
32'd28557: dataIn1 = 32'd35
; 
32'd28558: dataIn1 = 32'd38
; 
32'd28559: dataIn1 = 32'd39
; 
32'd28560: dataIn1 = 32'd42
; 
32'd28561: dataIn1 = 32'd44
; 
32'd28562: dataIn1 = 32'd45
; 
32'd28563: dataIn1 = 32'd46
; 
32'd28564: dataIn1 = 32'd47
; 
32'd28565: dataIn1 = 32'd48
; 
32'd28566: dataIn1 = 32'd53
; 
32'd28567: dataIn1 = 32'd54
; 
32'd28568: dataIn1 = 32'd55
; 
32'd28569: dataIn1 = 32'd56
; 
32'd28570: dataIn1 = 32'd57
; 
32'd28571: dataIn1 = 32'd58
; 
32'd28572: dataIn1 = 32'd59
; 
32'd28573: dataIn1 = 32'd60
; 
32'd28574: dataIn1 = 32'd61
; 
32'd28575: dataIn1 = 32'd0
; 
32'd28576: dataIn1 = 32'd1
; 
32'd28577: dataIn1 = 32'd3
; 
32'd28578: dataIn1 = 32'd4
; 
32'd28579: dataIn1 = 32'd5
; 
32'd28580: dataIn1 = 32'd6
; 
32'd28581: dataIn1 = 32'd12
; 
32'd28582: dataIn1 = 32'd13
; 
32'd28583: dataIn1 = 32'd14
; 
32'd28584: dataIn1 = 32'd15
; 
32'd28585: dataIn1 = 32'd16
; 
32'd28586: dataIn1 = 32'd19
; 
32'd28587: dataIn1 = 32'd20
; 
32'd28588: dataIn1 = 32'd23
; 
32'd28589: dataIn1 = 32'd24
; 
32'd28590: dataIn1 = 32'd28
; 
32'd28591: dataIn1 = 32'd30
; 
32'd28592: dataIn1 = 32'd31
; 
32'd28593: dataIn1 = 32'd32
; 
32'd28594: dataIn1 = 32'd34
; 
32'd28595: dataIn1 = 32'd35
; 
32'd28596: dataIn1 = 32'd37
; 
32'd28597: dataIn1 = 32'd38
; 
32'd28598: dataIn1 = 32'd39
; 
32'd28599: dataIn1 = 32'd40
; 
32'd28600: dataIn1 = 32'd41
; 
32'd28601: dataIn1 = 32'd42
; 
32'd28602: dataIn1 = 32'd43
; 
32'd28603: dataIn1 = 32'd45
; 
32'd28604: dataIn1 = 32'd46
; 
32'd28605: dataIn1 = 32'd49
; 
32'd28606: dataIn1 = 32'd50
; 
32'd28607: dataIn1 = 32'd55
; 
32'd28608: dataIn1 = 32'd58
; 
32'd28609: dataIn1 = 32'd60
; 
32'd28610: dataIn1 = 32'd61
; 
32'd28611: dataIn1 = 32'd62
; 
32'd28612: dataIn1 = 32'd63
; 
32'd28613: dataIn1 = 32'd1
; 
32'd28614: dataIn1 = 32'd4
; 
32'd28615: dataIn1 = 32'd5
; 
32'd28616: dataIn1 = 32'd6
; 
32'd28617: dataIn1 = 32'd8
; 
32'd28618: dataIn1 = 32'd12
; 
32'd28619: dataIn1 = 32'd13
; 
32'd28620: dataIn1 = 32'd14
; 
32'd28621: dataIn1 = 32'd16
; 
32'd28622: dataIn1 = 32'd17
; 
32'd28623: dataIn1 = 32'd18
; 
32'd28624: dataIn1 = 32'd19
; 
32'd28625: dataIn1 = 32'd21
; 
32'd28626: dataIn1 = 32'd23
; 
32'd28627: dataIn1 = 32'd28
; 
32'd28628: dataIn1 = 32'd29
; 
32'd28629: dataIn1 = 32'd31
; 
32'd28630: dataIn1 = 32'd32
; 
32'd28631: dataIn1 = 32'd33
; 
32'd28632: dataIn1 = 32'd34
; 
32'd28633: dataIn1 = 32'd35
; 
32'd28634: dataIn1 = 32'd39
; 
32'd28635: dataIn1 = 32'd40
; 
32'd28636: dataIn1 = 32'd43
; 
32'd28637: dataIn1 = 32'd44
; 
32'd28638: dataIn1 = 32'd46
; 
32'd28639: dataIn1 = 32'd47
; 
32'd28640: dataIn1 = 32'd48
; 
32'd28641: dataIn1 = 32'd49
; 
32'd28642: dataIn1 = 32'd52
; 
32'd28643: dataIn1 = 32'd53
; 
32'd28644: dataIn1 = 32'd55
; 
32'd28645: dataIn1 = 32'd56
; 
32'd28646: dataIn1 = 32'd57
; 
32'd28647: dataIn1 = 32'd61
; 
32'd28648: dataIn1 = 32'd62
; 
32'd28649: dataIn1 = 32'd63
; 
32'd28650: dataIn1 = 32'd1
; 
32'd28651: dataIn1 = 32'd2
; 
32'd28652: dataIn1 = 32'd4
; 
32'd28653: dataIn1 = 32'd6
; 
32'd28654: dataIn1 = 32'd10
; 
32'd28655: dataIn1 = 32'd11
; 
32'd28656: dataIn1 = 32'd14
; 
32'd28657: dataIn1 = 32'd15
; 
32'd28658: dataIn1 = 32'd16
; 
32'd28659: dataIn1 = 32'd19
; 
32'd28660: dataIn1 = 32'd20
; 
32'd28661: dataIn1 = 32'd21
; 
32'd28662: dataIn1 = 32'd22
; 
32'd28663: dataIn1 = 32'd23
; 
32'd28664: dataIn1 = 32'd24
; 
32'd28665: dataIn1 = 32'd25
; 
32'd28666: dataIn1 = 32'd26
; 
32'd28667: dataIn1 = 32'd27
; 
32'd28668: dataIn1 = 32'd28
; 
32'd28669: dataIn1 = 32'd29
; 
32'd28670: dataIn1 = 32'd31
; 
32'd28671: dataIn1 = 32'd33
; 
32'd28672: dataIn1 = 32'd34
; 
32'd28673: dataIn1 = 32'd35
; 
32'd28674: dataIn1 = 32'd36
; 
32'd28675: dataIn1 = 32'd37
; 
32'd28676: dataIn1 = 32'd38
; 
32'd28677: dataIn1 = 32'd41
; 
32'd28678: dataIn1 = 32'd43
; 
32'd28679: dataIn1 = 32'd44
; 
32'd28680: dataIn1 = 32'd45
; 
32'd28681: dataIn1 = 32'd46
; 
32'd28682: dataIn1 = 32'd49
; 
32'd28683: dataIn1 = 32'd51
; 
32'd28684: dataIn1 = 32'd52
; 
32'd28685: dataIn1 = 32'd55
; 
32'd28686: dataIn1 = 32'd58
; 
32'd28687: dataIn1 = 32'd60
; 
32'd28688: dataIn1 = 32'd62
; 
32'd28689: dataIn1 = 32'd63
; 
32'd28690: dataIn1 = 32'd1
; 
32'd28691: dataIn1 = 32'd3
; 
32'd28692: dataIn1 = 32'd4
; 
32'd28693: dataIn1 = 32'd7
; 
32'd28694: dataIn1 = 32'd10
; 
32'd28695: dataIn1 = 32'd12
; 
32'd28696: dataIn1 = 32'd13
; 
32'd28697: dataIn1 = 32'd14
; 
32'd28698: dataIn1 = 32'd15
; 
32'd28699: dataIn1 = 32'd16
; 
32'd28700: dataIn1 = 32'd19
; 
32'd28701: dataIn1 = 32'd20
; 
32'd28702: dataIn1 = 32'd21
; 
32'd28703: dataIn1 = 32'd23
; 
32'd28704: dataIn1 = 32'd24
; 
32'd28705: dataIn1 = 32'd26
; 
32'd28706: dataIn1 = 32'd28
; 
32'd28707: dataIn1 = 32'd29
; 
32'd28708: dataIn1 = 32'd30
; 
32'd28709: dataIn1 = 32'd31
; 
32'd28710: dataIn1 = 32'd33
; 
32'd28711: dataIn1 = 32'd35
; 
32'd28712: dataIn1 = 32'd39
; 
32'd28713: dataIn1 = 32'd41
; 
32'd28714: dataIn1 = 32'd43
; 
32'd28715: dataIn1 = 32'd44
; 
32'd28716: dataIn1 = 32'd48
; 
32'd28717: dataIn1 = 32'd50
; 
32'd28718: dataIn1 = 32'd52
; 
32'd28719: dataIn1 = 32'd55
; 
32'd28720: dataIn1 = 32'd56
; 
32'd28721: dataIn1 = 32'd59
; 
32'd28722: dataIn1 = 32'd60
; 
32'd28723: dataIn1 = 32'd61
; 
32'd28724: dataIn1 = 32'd62
; 
32'd28725: dataIn1 = 32'd1
; 
32'd28726: dataIn1 = 32'd2
; 
32'd28727: dataIn1 = 32'd3
; 
32'd28728: dataIn1 = 32'd4
; 
32'd28729: dataIn1 = 32'd5
; 
32'd28730: dataIn1 = 32'd7
; 
32'd28731: dataIn1 = 32'd11
; 
32'd28732: dataIn1 = 32'd12
; 
32'd28733: dataIn1 = 32'd15
; 
32'd28734: dataIn1 = 32'd16
; 
32'd28735: dataIn1 = 32'd18
; 
32'd28736: dataIn1 = 32'd20
; 
32'd28737: dataIn1 = 32'd21
; 
32'd28738: dataIn1 = 32'd23
; 
32'd28739: dataIn1 = 32'd24
; 
32'd28740: dataIn1 = 32'd25
; 
32'd28741: dataIn1 = 32'd28
; 
32'd28742: dataIn1 = 32'd29
; 
32'd28743: dataIn1 = 32'd33
; 
32'd28744: dataIn1 = 32'd35
; 
32'd28745: dataIn1 = 32'd40
; 
32'd28746: dataIn1 = 32'd44
; 
32'd28747: dataIn1 = 32'd47
; 
32'd28748: dataIn1 = 32'd48
; 
32'd28749: dataIn1 = 32'd49
; 
32'd28750: dataIn1 = 32'd51
; 
32'd28751: dataIn1 = 32'd56
; 
32'd28752: dataIn1 = 32'd57
; 
32'd28753: dataIn1 = 32'd58
; 
32'd28754: dataIn1 = 32'd59
; 
32'd28755: dataIn1 = 32'd1
; 
32'd28756: dataIn1 = 32'd4
; 
32'd28757: dataIn1 = 32'd5
; 
32'd28758: dataIn1 = 32'd6
; 
32'd28759: dataIn1 = 32'd7
; 
32'd28760: dataIn1 = 32'd9
; 
32'd28761: dataIn1 = 32'd13
; 
32'd28762: dataIn1 = 32'd16
; 
32'd28763: dataIn1 = 32'd17
; 
32'd28764: dataIn1 = 32'd18
; 
32'd28765: dataIn1 = 32'd21
; 
32'd28766: dataIn1 = 32'd23
; 
32'd28767: dataIn1 = 32'd24
; 
32'd28768: dataIn1 = 32'd26
; 
32'd28769: dataIn1 = 32'd27
; 
32'd28770: dataIn1 = 32'd30
; 
32'd28771: dataIn1 = 32'd32
; 
32'd28772: dataIn1 = 32'd33
; 
32'd28773: dataIn1 = 32'd35
; 
32'd28774: dataIn1 = 32'd36
; 
32'd28775: dataIn1 = 32'd38
; 
32'd28776: dataIn1 = 32'd39
; 
32'd28777: dataIn1 = 32'd40
; 
32'd28778: dataIn1 = 32'd42
; 
32'd28779: dataIn1 = 32'd43
; 
32'd28780: dataIn1 = 32'd46
; 
32'd28781: dataIn1 = 32'd49
; 
32'd28782: dataIn1 = 32'd53
; 
32'd28783: dataIn1 = 32'd55
; 
32'd28784: dataIn1 = 32'd57
; 
32'd28785: dataIn1 = 32'd58
; 
32'd28786: dataIn1 = 32'd59
; 
32'd28787: dataIn1 = 32'd62
; 
32'd28788: dataIn1 = 32'd63
; 
32'd28789: dataIn1 = 32'd0
; 
32'd28790: dataIn1 = 32'd1
; 
32'd28791: dataIn1 = 32'd2
; 
32'd28792: dataIn1 = 32'd6
; 
32'd28793: dataIn1 = 32'd7
; 
32'd28794: dataIn1 = 32'd9
; 
32'd28795: dataIn1 = 32'd10
; 
32'd28796: dataIn1 = 32'd11
; 
32'd28797: dataIn1 = 32'd14
; 
32'd28798: dataIn1 = 32'd15
; 
32'd28799: dataIn1 = 32'd20
; 
32'd28800: dataIn1 = 32'd23
; 
32'd28801: dataIn1 = 32'd24
; 
32'd28802: dataIn1 = 32'd25
; 
32'd28803: dataIn1 = 32'd27
; 
32'd28804: dataIn1 = 32'd28
; 
32'd28805: dataIn1 = 32'd31
; 
32'd28806: dataIn1 = 32'd33
; 
32'd28807: dataIn1 = 32'd34
; 
32'd28808: dataIn1 = 32'd36
; 
32'd28809: dataIn1 = 32'd39
; 
32'd28810: dataIn1 = 32'd41
; 
32'd28811: dataIn1 = 32'd42
; 
32'd28812: dataIn1 = 32'd44
; 
32'd28813: dataIn1 = 32'd45
; 
32'd28814: dataIn1 = 32'd46
; 
32'd28815: dataIn1 = 32'd47
; 
32'd28816: dataIn1 = 32'd48
; 
32'd28817: dataIn1 = 32'd55
; 
32'd28818: dataIn1 = 32'd56
; 
32'd28819: dataIn1 = 32'd57
; 
32'd28820: dataIn1 = 32'd58
; 
32'd28821: dataIn1 = 32'd62
; 
32'd28822: dataIn1 = 32'd63
; 
32'd28823: dataIn1 = 32'd2
; 
32'd28824: dataIn1 = 32'd3
; 
32'd28825: dataIn1 = 32'd5
; 
32'd28826: dataIn1 = 32'd7
; 
32'd28827: dataIn1 = 32'd8
; 
32'd28828: dataIn1 = 32'd11
; 
32'd28829: dataIn1 = 32'd12
; 
32'd28830: dataIn1 = 32'd13
; 
32'd28831: dataIn1 = 32'd14
; 
32'd28832: dataIn1 = 32'd17
; 
32'd28833: dataIn1 = 32'd18
; 
32'd28834: dataIn1 = 32'd20
; 
32'd28835: dataIn1 = 32'd21
; 
32'd28836: dataIn1 = 32'd22
; 
32'd28837: dataIn1 = 32'd23
; 
32'd28838: dataIn1 = 32'd29
; 
32'd28839: dataIn1 = 32'd30
; 
32'd28840: dataIn1 = 32'd32
; 
32'd28841: dataIn1 = 32'd33
; 
32'd28842: dataIn1 = 32'd36
; 
32'd28843: dataIn1 = 32'd38
; 
32'd28844: dataIn1 = 32'd39
; 
32'd28845: dataIn1 = 32'd43
; 
32'd28846: dataIn1 = 32'd44
; 
32'd28847: dataIn1 = 32'd45
; 
32'd28848: dataIn1 = 32'd46
; 
32'd28849: dataIn1 = 32'd47
; 
32'd28850: dataIn1 = 32'd49
; 
32'd28851: dataIn1 = 32'd51
; 
32'd28852: dataIn1 = 32'd53
; 
32'd28853: dataIn1 = 32'd56
; 
32'd28854: dataIn1 = 32'd57
; 
32'd28855: dataIn1 = 32'd62
; 
32'd28856: dataIn1 = 32'd63
; 
32'd28857: dataIn1 = 32'd2
; 
32'd28858: dataIn1 = 32'd3
; 
32'd28859: dataIn1 = 32'd6
; 
32'd28860: dataIn1 = 32'd8
; 
32'd28861: dataIn1 = 32'd10
; 
32'd28862: dataIn1 = 32'd11
; 
32'd28863: dataIn1 = 32'd14
; 
32'd28864: dataIn1 = 32'd16
; 
32'd28865: dataIn1 = 32'd19
; 
32'd28866: dataIn1 = 32'd23
; 
32'd28867: dataIn1 = 32'd24
; 
32'd28868: dataIn1 = 32'd26
; 
32'd28869: dataIn1 = 32'd27
; 
32'd28870: dataIn1 = 32'd32
; 
32'd28871: dataIn1 = 32'd34
; 
32'd28872: dataIn1 = 32'd36
; 
32'd28873: dataIn1 = 32'd38
; 
32'd28874: dataIn1 = 32'd39
; 
32'd28875: dataIn1 = 32'd40
; 
32'd28876: dataIn1 = 32'd42
; 
32'd28877: dataIn1 = 32'd43
; 
32'd28878: dataIn1 = 32'd44
; 
32'd28879: dataIn1 = 32'd46
; 
32'd28880: dataIn1 = 32'd47
; 
32'd28881: dataIn1 = 32'd49
; 
32'd28882: dataIn1 = 32'd51
; 
32'd28883: dataIn1 = 32'd57
; 
32'd28884: dataIn1 = 32'd58
; 
32'd28885: dataIn1 = 32'd59
; 
32'd28886: dataIn1 = 32'd62
; 
32'd28887: dataIn1 = 32'd0
; 
32'd28888: dataIn1 = 32'd2
; 
32'd28889: dataIn1 = 32'd3
; 
32'd28890: dataIn1 = 32'd5
; 
32'd28891: dataIn1 = 32'd6
; 
32'd28892: dataIn1 = 32'd7
; 
32'd28893: dataIn1 = 32'd8
; 
32'd28894: dataIn1 = 32'd9
; 
32'd28895: dataIn1 = 32'd12
; 
32'd28896: dataIn1 = 32'd13
; 
32'd28897: dataIn1 = 32'd14
; 
32'd28898: dataIn1 = 32'd15
; 
32'd28899: dataIn1 = 32'd16
; 
32'd28900: dataIn1 = 32'd18
; 
32'd28901: dataIn1 = 32'd19
; 
32'd28902: dataIn1 = 32'd21
; 
32'd28903: dataIn1 = 32'd26
; 
32'd28904: dataIn1 = 32'd27
; 
32'd28905: dataIn1 = 32'd34
; 
32'd28906: dataIn1 = 32'd35
; 
32'd28907: dataIn1 = 32'd40
; 
32'd28908: dataIn1 = 32'd42
; 
32'd28909: dataIn1 = 32'd44
; 
32'd28910: dataIn1 = 32'd45
; 
32'd28911: dataIn1 = 32'd46
; 
32'd28912: dataIn1 = 32'd47
; 
32'd28913: dataIn1 = 32'd48
; 
32'd28914: dataIn1 = 32'd49
; 
32'd28915: dataIn1 = 32'd50
; 
32'd28916: dataIn1 = 32'd51
; 
32'd28917: dataIn1 = 32'd52
; 
32'd28918: dataIn1 = 32'd54
; 
32'd28919: dataIn1 = 32'd55
; 
32'd28920: dataIn1 = 32'd56
; 
32'd28921: dataIn1 = 32'd57
; 
32'd28922: dataIn1 = 32'd58
; 
32'd28923: dataIn1 = 32'd59
; 
32'd28924: dataIn1 = 32'd60
; 
32'd28925: dataIn1 = 32'd61
; 
32'd28926: dataIn1 = 32'd62
; 
32'd28927: dataIn1 = 32'd63
; 
32'd28928: dataIn1 = 32'd0
; 
32'd28929: dataIn1 = 32'd2
; 
32'd28930: dataIn1 = 32'd3
; 
32'd28931: dataIn1 = 32'd6
; 
32'd28932: dataIn1 = 32'd7
; 
32'd28933: dataIn1 = 32'd8
; 
32'd28934: dataIn1 = 32'd9
; 
32'd28935: dataIn1 = 32'd10
; 
32'd28936: dataIn1 = 32'd12
; 
32'd28937: dataIn1 = 32'd13
; 
32'd28938: dataIn1 = 32'd14
; 
32'd28939: dataIn1 = 32'd15
; 
32'd28940: dataIn1 = 32'd20
; 
32'd28941: dataIn1 = 32'd23
; 
32'd28942: dataIn1 = 32'd24
; 
32'd28943: dataIn1 = 32'd30
; 
32'd28944: dataIn1 = 32'd33
; 
32'd28945: dataIn1 = 32'd34
; 
32'd28946: dataIn1 = 32'd36
; 
32'd28947: dataIn1 = 32'd37
; 
32'd28948: dataIn1 = 32'd40
; 
32'd28949: dataIn1 = 32'd41
; 
32'd28950: dataIn1 = 32'd43
; 
32'd28951: dataIn1 = 32'd45
; 
32'd28952: dataIn1 = 32'd47
; 
32'd28953: dataIn1 = 32'd48
; 
32'd28954: dataIn1 = 32'd49
; 
32'd28955: dataIn1 = 32'd50
; 
32'd28956: dataIn1 = 32'd51
; 
32'd28957: dataIn1 = 32'd54
; 
32'd28958: dataIn1 = 32'd57
; 
32'd28959: dataIn1 = 32'd58
; 
32'd28960: dataIn1 = 32'd59
; 
32'd28961: dataIn1 = 32'd60
; 
32'd28962: dataIn1 = 32'd61
; 
32'd28963: dataIn1 = 32'd0
; 
32'd28964: dataIn1 = 32'd1
; 
32'd28965: dataIn1 = 32'd3
; 
32'd28966: dataIn1 = 32'd4
; 
32'd28967: dataIn1 = 32'd5
; 
32'd28968: dataIn1 = 32'd6
; 
32'd28969: dataIn1 = 32'd8
; 
32'd28970: dataIn1 = 32'd9
; 
32'd28971: dataIn1 = 32'd10
; 
32'd28972: dataIn1 = 32'd11
; 
32'd28973: dataIn1 = 32'd13
; 
32'd28974: dataIn1 = 32'd19
; 
32'd28975: dataIn1 = 32'd20
; 
32'd28976: dataIn1 = 32'd21
; 
32'd28977: dataIn1 = 32'd22
; 
32'd28978: dataIn1 = 32'd23
; 
32'd28979: dataIn1 = 32'd25
; 
32'd28980: dataIn1 = 32'd27
; 
32'd28981: dataIn1 = 32'd28
; 
32'd28982: dataIn1 = 32'd29
; 
32'd28983: dataIn1 = 32'd32
; 
32'd28984: dataIn1 = 32'd33
; 
32'd28985: dataIn1 = 32'd34
; 
32'd28986: dataIn1 = 32'd35
; 
32'd28987: dataIn1 = 32'd36
; 
32'd28988: dataIn1 = 32'd38
; 
32'd28989: dataIn1 = 32'd39
; 
32'd28990: dataIn1 = 32'd42
; 
32'd28991: dataIn1 = 32'd43
; 
32'd28992: dataIn1 = 32'd44
; 
32'd28993: dataIn1 = 32'd45
; 
32'd28994: dataIn1 = 32'd46
; 
32'd28995: dataIn1 = 32'd48
; 
32'd28996: dataIn1 = 32'd49
; 
32'd28997: dataIn1 = 32'd51
; 
32'd28998: dataIn1 = 32'd52
; 
32'd28999: dataIn1 = 32'd53
; 
32'd29000: dataIn1 = 32'd55
; 
32'd29001: dataIn1 = 32'd56
; 
32'd29002: dataIn1 = 32'd57
; 
32'd29003: dataIn1 = 32'd60
; 
32'd29004: dataIn1 = 32'd61
; 
32'd29005: dataIn1 = 32'd62
; 
32'd29006: dataIn1 = 32'd63
; 
32'd29007: dataIn1 = 32'd0
; 
32'd29008: dataIn1 = 32'd1
; 
32'd29009: dataIn1 = 32'd2
; 
32'd29010: dataIn1 = 32'd3
; 
32'd29011: dataIn1 = 32'd6
; 
32'd29012: dataIn1 = 32'd12
; 
32'd29013: dataIn1 = 32'd13
; 
32'd29014: dataIn1 = 32'd15
; 
32'd29015: dataIn1 = 32'd16
; 
32'd29016: dataIn1 = 32'd18
; 
32'd29017: dataIn1 = 32'd19
; 
32'd29018: dataIn1 = 32'd20
; 
32'd29019: dataIn1 = 32'd21
; 
32'd29020: dataIn1 = 32'd25
; 
32'd29021: dataIn1 = 32'd26
; 
32'd29022: dataIn1 = 32'd27
; 
32'd29023: dataIn1 = 32'd28
; 
32'd29024: dataIn1 = 32'd29
; 
32'd29025: dataIn1 = 32'd30
; 
32'd29026: dataIn1 = 32'd31
; 
32'd29027: dataIn1 = 32'd33
; 
32'd29028: dataIn1 = 32'd34
; 
32'd29029: dataIn1 = 32'd37
; 
32'd29030: dataIn1 = 32'd38
; 
32'd29031: dataIn1 = 32'd40
; 
32'd29032: dataIn1 = 32'd42
; 
32'd29033: dataIn1 = 32'd45
; 
32'd29034: dataIn1 = 32'd46
; 
32'd29035: dataIn1 = 32'd48
; 
32'd29036: dataIn1 = 32'd50
; 
32'd29037: dataIn1 = 32'd52
; 
32'd29038: dataIn1 = 32'd54
; 
32'd29039: dataIn1 = 32'd55
; 
32'd29040: dataIn1 = 32'd59
; 
32'd29041: dataIn1 = 32'd60
; 
32'd29042: dataIn1 = 32'd63
; 
32'd29043: dataIn1 = 32'd0
; 
32'd29044: dataIn1 = 32'd1
; 
32'd29045: dataIn1 = 32'd2
; 
32'd29046: dataIn1 = 32'd4
; 
32'd29047: dataIn1 = 32'd5
; 
32'd29048: dataIn1 = 32'd7
; 
32'd29049: dataIn1 = 32'd8
; 
32'd29050: dataIn1 = 32'd9
; 
32'd29051: dataIn1 = 32'd11
; 
32'd29052: dataIn1 = 32'd15
; 
32'd29053: dataIn1 = 32'd16
; 
32'd29054: dataIn1 = 32'd18
; 
32'd29055: dataIn1 = 32'd23
; 
32'd29056: dataIn1 = 32'd25
; 
32'd29057: dataIn1 = 32'd27
; 
32'd29058: dataIn1 = 32'd30
; 
32'd29059: dataIn1 = 32'd31
; 
32'd29060: dataIn1 = 32'd32
; 
32'd29061: dataIn1 = 32'd33
; 
32'd29062: dataIn1 = 32'd37
; 
32'd29063: dataIn1 = 32'd42
; 
32'd29064: dataIn1 = 32'd45
; 
32'd29065: dataIn1 = 32'd46
; 
32'd29066: dataIn1 = 32'd49
; 
32'd29067: dataIn1 = 32'd51
; 
32'd29068: dataIn1 = 32'd52
; 
32'd29069: dataIn1 = 32'd53
; 
32'd29070: dataIn1 = 32'd54
; 
32'd29071: dataIn1 = 32'd55
; 
32'd29072: dataIn1 = 32'd56
; 
32'd29073: dataIn1 = 32'd59
; 
32'd29074: dataIn1 = 32'd63
; 
32'd29075: dataIn1 = 32'd0
; 
32'd29076: dataIn1 = 32'd1
; 
32'd29077: dataIn1 = 32'd3
; 
32'd29078: dataIn1 = 32'd5
; 
32'd29079: dataIn1 = 32'd6
; 
32'd29080: dataIn1 = 32'd7
; 
32'd29081: dataIn1 = 32'd8
; 
32'd29082: dataIn1 = 32'd10
; 
32'd29083: dataIn1 = 32'd11
; 
32'd29084: dataIn1 = 32'd12
; 
32'd29085: dataIn1 = 32'd14
; 
32'd29086: dataIn1 = 32'd15
; 
32'd29087: dataIn1 = 32'd17
; 
32'd29088: dataIn1 = 32'd18
; 
32'd29089: dataIn1 = 32'd21
; 
32'd29090: dataIn1 = 32'd23
; 
32'd29091: dataIn1 = 32'd24
; 
32'd29092: dataIn1 = 32'd25
; 
32'd29093: dataIn1 = 32'd26
; 
32'd29094: dataIn1 = 32'd28
; 
32'd29095: dataIn1 = 32'd30
; 
32'd29096: dataIn1 = 32'd31
; 
32'd29097: dataIn1 = 32'd32
; 
32'd29098: dataIn1 = 32'd33
; 
32'd29099: dataIn1 = 32'd35
; 
32'd29100: dataIn1 = 32'd37
; 
32'd29101: dataIn1 = 32'd39
; 
32'd29102: dataIn1 = 32'd40
; 
32'd29103: dataIn1 = 32'd41
; 
32'd29104: dataIn1 = 32'd42
; 
32'd29105: dataIn1 = 32'd43
; 
32'd29106: dataIn1 = 32'd48
; 
32'd29107: dataIn1 = 32'd49
; 
32'd29108: dataIn1 = 32'd50
; 
32'd29109: dataIn1 = 32'd51
; 
32'd29110: dataIn1 = 32'd54
; 
32'd29111: dataIn1 = 32'd56
; 
32'd29112: dataIn1 = 32'd57
; 
32'd29113: dataIn1 = 32'd58
; 
32'd29114: dataIn1 = 32'd60
; 
32'd29115: dataIn1 = 32'd62
; 
32'd29116: dataIn1 = 32'd63
; 
32'd29117: dataIn1 = 32'd4
; 
32'd29118: dataIn1 = 32'd6
; 
32'd29119: dataIn1 = 32'd8
; 
32'd29120: dataIn1 = 32'd10
; 
32'd29121: dataIn1 = 32'd12
; 
32'd29122: dataIn1 = 32'd14
; 
32'd29123: dataIn1 = 32'd15
; 
32'd29124: dataIn1 = 32'd19
; 
32'd29125: dataIn1 = 32'd20
; 
32'd29126: dataIn1 = 32'd21
; 
32'd29127: dataIn1 = 32'd22
; 
32'd29128: dataIn1 = 32'd23
; 
32'd29129: dataIn1 = 32'd24
; 
32'd29130: dataIn1 = 32'd25
; 
32'd29131: dataIn1 = 32'd26
; 
32'd29132: dataIn1 = 32'd27
; 
32'd29133: dataIn1 = 32'd28
; 
32'd29134: dataIn1 = 32'd31
; 
32'd29135: dataIn1 = 32'd32
; 
32'd29136: dataIn1 = 32'd33
; 
32'd29137: dataIn1 = 32'd35
; 
32'd29138: dataIn1 = 32'd36
; 
32'd29139: dataIn1 = 32'd40
; 
32'd29140: dataIn1 = 32'd43
; 
32'd29141: dataIn1 = 32'd44
; 
32'd29142: dataIn1 = 32'd45
; 
32'd29143: dataIn1 = 32'd48
; 
32'd29144: dataIn1 = 32'd51
; 
32'd29145: dataIn1 = 32'd52
; 
32'd29146: dataIn1 = 32'd54
; 
32'd29147: dataIn1 = 32'd55
; 
32'd29148: dataIn1 = 32'd56
; 
32'd29149: dataIn1 = 32'd58
; 
32'd29150: dataIn1 = 32'd60
; 
32'd29151: dataIn1 = 32'd61
; 
32'd29152: dataIn1 = 32'd62
; 
32'd29153: dataIn1 = 32'd63
; 
32'd29154: dataIn1 = 32'd2
; 
32'd29155: dataIn1 = 32'd4
; 
32'd29156: dataIn1 = 32'd5
; 
32'd29157: dataIn1 = 32'd7
; 
32'd29158: dataIn1 = 32'd8
; 
32'd29159: dataIn1 = 32'd10
; 
32'd29160: dataIn1 = 32'd11
; 
32'd29161: dataIn1 = 32'd12
; 
32'd29162: dataIn1 = 32'd15
; 
32'd29163: dataIn1 = 32'd16
; 
32'd29164: dataIn1 = 32'd17
; 
32'd29165: dataIn1 = 32'd19
; 
32'd29166: dataIn1 = 32'd23
; 
32'd29167: dataIn1 = 32'd24
; 
32'd29168: dataIn1 = 32'd25
; 
32'd29169: dataIn1 = 32'd26
; 
32'd29170: dataIn1 = 32'd27
; 
32'd29171: dataIn1 = 32'd29
; 
32'd29172: dataIn1 = 32'd31
; 
32'd29173: dataIn1 = 32'd32
; 
32'd29174: dataIn1 = 32'd34
; 
32'd29175: dataIn1 = 32'd36
; 
32'd29176: dataIn1 = 32'd38
; 
32'd29177: dataIn1 = 32'd40
; 
32'd29178: dataIn1 = 32'd42
; 
32'd29179: dataIn1 = 32'd43
; 
32'd29180: dataIn1 = 32'd46
; 
32'd29181: dataIn1 = 32'd47
; 
32'd29182: dataIn1 = 32'd49
; 
32'd29183: dataIn1 = 32'd51
; 
32'd29184: dataIn1 = 32'd52
; 
32'd29185: dataIn1 = 32'd53
; 
32'd29186: dataIn1 = 32'd54
; 
32'd29187: dataIn1 = 32'd55
; 
32'd29188: dataIn1 = 32'd57
; 
32'd29189: dataIn1 = 32'd58
; 
32'd29190: dataIn1 = 32'd61
; 
32'd29191: dataIn1 = 32'd62
; 
32'd29192: dataIn1 = 32'd63
; 
32'd29193: dataIn1 = 32'd0
; 
32'd29194: dataIn1 = 32'd1
; 
32'd29195: dataIn1 = 32'd2
; 
32'd29196: dataIn1 = 32'd3
; 
32'd29197: dataIn1 = 32'd5
; 
32'd29198: dataIn1 = 32'd11
; 
32'd29199: dataIn1 = 32'd13
; 
32'd29200: dataIn1 = 32'd14
; 
32'd29201: dataIn1 = 32'd15
; 
32'd29202: dataIn1 = 32'd17
; 
32'd29203: dataIn1 = 32'd19
; 
32'd29204: dataIn1 = 32'd23
; 
32'd29205: dataIn1 = 32'd27
; 
32'd29206: dataIn1 = 32'd29
; 
32'd29207: dataIn1 = 32'd30
; 
32'd29208: dataIn1 = 32'd32
; 
32'd29209: dataIn1 = 32'd33
; 
32'd29210: dataIn1 = 32'd35
; 
32'd29211: dataIn1 = 32'd36
; 
32'd29212: dataIn1 = 32'd37
; 
32'd29213: dataIn1 = 32'd38
; 
32'd29214: dataIn1 = 32'd39
; 
32'd29215: dataIn1 = 32'd41
; 
32'd29216: dataIn1 = 32'd48
; 
32'd29217: dataIn1 = 32'd50
; 
32'd29218: dataIn1 = 32'd51
; 
32'd29219: dataIn1 = 32'd52
; 
32'd29220: dataIn1 = 32'd53
; 
32'd29221: dataIn1 = 32'd54
; 
32'd29222: dataIn1 = 32'd55
; 
32'd29223: dataIn1 = 32'd56
; 
32'd29224: dataIn1 = 32'd58
; 
32'd29225: dataIn1 = 32'd60
; 
32'd29226: dataIn1 = 32'd62
; 
32'd29227: dataIn1 = 32'd0
; 
32'd29228: dataIn1 = 32'd1
; 
32'd29229: dataIn1 = 32'd2
; 
32'd29230: dataIn1 = 32'd3
; 
32'd29231: dataIn1 = 32'd5
; 
32'd29232: dataIn1 = 32'd9
; 
32'd29233: dataIn1 = 32'd13
; 
32'd29234: dataIn1 = 32'd14
; 
32'd29235: dataIn1 = 32'd15
; 
32'd29236: dataIn1 = 32'd16
; 
32'd29237: dataIn1 = 32'd18
; 
32'd29238: dataIn1 = 32'd19
; 
32'd29239: dataIn1 = 32'd20
; 
32'd29240: dataIn1 = 32'd21
; 
32'd29241: dataIn1 = 32'd22
; 
32'd29242: dataIn1 = 32'd24
; 
32'd29243: dataIn1 = 32'd26
; 
32'd29244: dataIn1 = 32'd31
; 
32'd29245: dataIn1 = 32'd33
; 
32'd29246: dataIn1 = 32'd34
; 
32'd29247: dataIn1 = 32'd36
; 
32'd29248: dataIn1 = 32'd37
; 
32'd29249: dataIn1 = 32'd42
; 
32'd29250: dataIn1 = 32'd43
; 
32'd29251: dataIn1 = 32'd45
; 
32'd29252: dataIn1 = 32'd46
; 
32'd29253: dataIn1 = 32'd47
; 
32'd29254: dataIn1 = 32'd49
; 
32'd29255: dataIn1 = 32'd51
; 
32'd29256: dataIn1 = 32'd56
; 
32'd29257: dataIn1 = 32'd57
; 
32'd29258: dataIn1 = 32'd58
; 
32'd29259: dataIn1 = 32'd62
; 
32'd29260: dataIn1 = 32'd0
; 
32'd29261: dataIn1 = 32'd1
; 
32'd29262: dataIn1 = 32'd2
; 
32'd29263: dataIn1 = 32'd3
; 
32'd29264: dataIn1 = 32'd4
; 
32'd29265: dataIn1 = 32'd5
; 
32'd29266: dataIn1 = 32'd7
; 
32'd29267: dataIn1 = 32'd8
; 
32'd29268: dataIn1 = 32'd10
; 
32'd29269: dataIn1 = 32'd14
; 
32'd29270: dataIn1 = 32'd15
; 
32'd29271: dataIn1 = 32'd20
; 
32'd29272: dataIn1 = 32'd21
; 
32'd29273: dataIn1 = 32'd24
; 
32'd29274: dataIn1 = 32'd25
; 
32'd29275: dataIn1 = 32'd27
; 
32'd29276: dataIn1 = 32'd28
; 
32'd29277: dataIn1 = 32'd29
; 
32'd29278: dataIn1 = 32'd32
; 
32'd29279: dataIn1 = 32'd33
; 
32'd29280: dataIn1 = 32'd34
; 
32'd29281: dataIn1 = 32'd35
; 
32'd29282: dataIn1 = 32'd36
; 
32'd29283: dataIn1 = 32'd37
; 
32'd29284: dataIn1 = 32'd38
; 
32'd29285: dataIn1 = 32'd41
; 
32'd29286: dataIn1 = 32'd43
; 
32'd29287: dataIn1 = 32'd44
; 
32'd29288: dataIn1 = 32'd45
; 
32'd29289: dataIn1 = 32'd46
; 
32'd29290: dataIn1 = 32'd47
; 
32'd29291: dataIn1 = 32'd50
; 
32'd29292: dataIn1 = 32'd51
; 
32'd29293: dataIn1 = 32'd53
; 
32'd29294: dataIn1 = 32'd54
; 
32'd29295: dataIn1 = 32'd55
; 
32'd29296: dataIn1 = 32'd56
; 
32'd29297: dataIn1 = 32'd57
; 
32'd29298: dataIn1 = 32'd58
; 
32'd29299: dataIn1 = 32'd59
; 
32'd29300: dataIn1 = 32'd60
; 
32'd29301: dataIn1 = 32'd61
; 
32'd29302: dataIn1 = 32'd62
; 
32'd29303: dataIn1 = 32'd63
; 
32'd29304: dataIn1 = 32'd0
; 
32'd29305: dataIn1 = 32'd1
; 
32'd29306: dataIn1 = 32'd2
; 
32'd29307: dataIn1 = 32'd4
; 
32'd29308: dataIn1 = 32'd5
; 
32'd29309: dataIn1 = 32'd8
; 
32'd29310: dataIn1 = 32'd9
; 
32'd29311: dataIn1 = 32'd11
; 
32'd29312: dataIn1 = 32'd13
; 
32'd29313: dataIn1 = 32'd14
; 
32'd29314: dataIn1 = 32'd16
; 
32'd29315: dataIn1 = 32'd22
; 
32'd29316: dataIn1 = 32'd23
; 
32'd29317: dataIn1 = 32'd24
; 
32'd29318: dataIn1 = 32'd25
; 
32'd29319: dataIn1 = 32'd28
; 
32'd29320: dataIn1 = 32'd30
; 
32'd29321: dataIn1 = 32'd31
; 
32'd29322: dataIn1 = 32'd32
; 
32'd29323: dataIn1 = 32'd34
; 
32'd29324: dataIn1 = 32'd37
; 
32'd29325: dataIn1 = 32'd38
; 
32'd29326: dataIn1 = 32'd40
; 
32'd29327: dataIn1 = 32'd43
; 
32'd29328: dataIn1 = 32'd44
; 
32'd29329: dataIn1 = 32'd46
; 
32'd29330: dataIn1 = 32'd48
; 
32'd29331: dataIn1 = 32'd49
; 
32'd29332: dataIn1 = 32'd50
; 
32'd29333: dataIn1 = 32'd51
; 
32'd29334: dataIn1 = 32'd52
; 
32'd29335: dataIn1 = 32'd53
; 
32'd29336: dataIn1 = 32'd54
; 
32'd29337: dataIn1 = 32'd58
; 
32'd29338: dataIn1 = 32'd59
; 
32'd29339: dataIn1 = 32'd61
; 
32'd29340: dataIn1 = 32'd62
; 
32'd29341: dataIn1 = 32'd1
; 
32'd29342: dataIn1 = 32'd2
; 
32'd29343: dataIn1 = 32'd4
; 
32'd29344: dataIn1 = 32'd11
; 
32'd29345: dataIn1 = 32'd12
; 
32'd29346: dataIn1 = 32'd13
; 
32'd29347: dataIn1 = 32'd14
; 
32'd29348: dataIn1 = 32'd16
; 
32'd29349: dataIn1 = 32'd18
; 
32'd29350: dataIn1 = 32'd21
; 
32'd29351: dataIn1 = 32'd22
; 
32'd29352: dataIn1 = 32'd23
; 
32'd29353: dataIn1 = 32'd25
; 
32'd29354: dataIn1 = 32'd26
; 
32'd29355: dataIn1 = 32'd27
; 
32'd29356: dataIn1 = 32'd28
; 
32'd29357: dataIn1 = 32'd30
; 
32'd29358: dataIn1 = 32'd31
; 
32'd29359: dataIn1 = 32'd39
; 
32'd29360: dataIn1 = 32'd40
; 
32'd29361: dataIn1 = 32'd41
; 
32'd29362: dataIn1 = 32'd42
; 
32'd29363: dataIn1 = 32'd43
; 
32'd29364: dataIn1 = 32'd44
; 
32'd29365: dataIn1 = 32'd46
; 
32'd29366: dataIn1 = 32'd47
; 
32'd29367: dataIn1 = 32'd51
; 
32'd29368: dataIn1 = 32'd52
; 
32'd29369: dataIn1 = 32'd54
; 
32'd29370: dataIn1 = 32'd57
; 
32'd29371: dataIn1 = 32'd60
; 
32'd29372: dataIn1 = 32'd0
; 
32'd29373: dataIn1 = 32'd2
; 
32'd29374: dataIn1 = 32'd3
; 
32'd29375: dataIn1 = 32'd5
; 
32'd29376: dataIn1 = 32'd6
; 
32'd29377: dataIn1 = 32'd8
; 
32'd29378: dataIn1 = 32'd9
; 
32'd29379: dataIn1 = 32'd11
; 
32'd29380: dataIn1 = 32'd12
; 
32'd29381: dataIn1 = 32'd13
; 
32'd29382: dataIn1 = 32'd14
; 
32'd29383: dataIn1 = 32'd20
; 
32'd29384: dataIn1 = 32'd21
; 
32'd29385: dataIn1 = 32'd25
; 
32'd29386: dataIn1 = 32'd26
; 
32'd29387: dataIn1 = 32'd27
; 
32'd29388: dataIn1 = 32'd28
; 
32'd29389: dataIn1 = 32'd31
; 
32'd29390: dataIn1 = 32'd33
; 
32'd29391: dataIn1 = 32'd36
; 
32'd29392: dataIn1 = 32'd37
; 
32'd29393: dataIn1 = 32'd38
; 
32'd29394: dataIn1 = 32'd40
; 
32'd29395: dataIn1 = 32'd42
; 
32'd29396: dataIn1 = 32'd46
; 
32'd29397: dataIn1 = 32'd47
; 
32'd29398: dataIn1 = 32'd52
; 
32'd29399: dataIn1 = 32'd53
; 
32'd29400: dataIn1 = 32'd54
; 
32'd29401: dataIn1 = 32'd57
; 
32'd29402: dataIn1 = 32'd58
; 
32'd29403: dataIn1 = 32'd59
; 
32'd29404: dataIn1 = 32'd61
; 
32'd29405: dataIn1 = 32'd0
; 
32'd29406: dataIn1 = 32'd2
; 
32'd29407: dataIn1 = 32'd3
; 
32'd29408: dataIn1 = 32'd5
; 
32'd29409: dataIn1 = 32'd7
; 
32'd29410: dataIn1 = 32'd9
; 
32'd29411: dataIn1 = 32'd14
; 
32'd29412: dataIn1 = 32'd16
; 
32'd29413: dataIn1 = 32'd17
; 
32'd29414: dataIn1 = 32'd18
; 
32'd29415: dataIn1 = 32'd20
; 
32'd29416: dataIn1 = 32'd21
; 
32'd29417: dataIn1 = 32'd22
; 
32'd29418: dataIn1 = 32'd24
; 
32'd29419: dataIn1 = 32'd25
; 
32'd29420: dataIn1 = 32'd27
; 
32'd29421: dataIn1 = 32'd29
; 
32'd29422: dataIn1 = 32'd30
; 
32'd29423: dataIn1 = 32'd33
; 
32'd29424: dataIn1 = 32'd34
; 
32'd29425: dataIn1 = 32'd36
; 
32'd29426: dataIn1 = 32'd37
; 
32'd29427: dataIn1 = 32'd41
; 
32'd29428: dataIn1 = 32'd42
; 
32'd29429: dataIn1 = 32'd45
; 
32'd29430: dataIn1 = 32'd46
; 
32'd29431: dataIn1 = 32'd47
; 
32'd29432: dataIn1 = 32'd49
; 
32'd29433: dataIn1 = 32'd50
; 
32'd29434: dataIn1 = 32'd52
; 
32'd29435: dataIn1 = 32'd53
; 
32'd29436: dataIn1 = 32'd54
; 
32'd29437: dataIn1 = 32'd55
; 
32'd29438: dataIn1 = 32'd57
; 
32'd29439: dataIn1 = 32'd58
; 
32'd29440: dataIn1 = 32'd60
; 
32'd29441: dataIn1 = 32'd61
; 
32'd29442: dataIn1 = 32'd63
; 
32'd29443: dataIn1 = 32'd0
; 
32'd29444: dataIn1 = 32'd1
; 
32'd29445: dataIn1 = 32'd2
; 
32'd29446: dataIn1 = 32'd5
; 
32'd29447: dataIn1 = 32'd8
; 
32'd29448: dataIn1 = 32'd11
; 
32'd29449: dataIn1 = 32'd12
; 
32'd29450: dataIn1 = 32'd13
; 
32'd29451: dataIn1 = 32'd15
; 
32'd29452: dataIn1 = 32'd17
; 
32'd29453: dataIn1 = 32'd18
; 
32'd29454: dataIn1 = 32'd20
; 
32'd29455: dataIn1 = 32'd21
; 
32'd29456: dataIn1 = 32'd22
; 
32'd29457: dataIn1 = 32'd24
; 
32'd29458: dataIn1 = 32'd25
; 
32'd29459: dataIn1 = 32'd26
; 
32'd29460: dataIn1 = 32'd28
; 
32'd29461: dataIn1 = 32'd29
; 
32'd29462: dataIn1 = 32'd30
; 
32'd29463: dataIn1 = 32'd34
; 
32'd29464: dataIn1 = 32'd35
; 
32'd29465: dataIn1 = 32'd38
; 
32'd29466: dataIn1 = 32'd39
; 
32'd29467: dataIn1 = 32'd41
; 
32'd29468: dataIn1 = 32'd43
; 
32'd29469: dataIn1 = 32'd45
; 
32'd29470: dataIn1 = 32'd46
; 
32'd29471: dataIn1 = 32'd48
; 
32'd29472: dataIn1 = 32'd50
; 
32'd29473: dataIn1 = 32'd51
; 
32'd29474: dataIn1 = 32'd52
; 
32'd29475: dataIn1 = 32'd53
; 
32'd29476: dataIn1 = 32'd54
; 
32'd29477: dataIn1 = 32'd56
; 
32'd29478: dataIn1 = 32'd58
; 
32'd29479: dataIn1 = 32'd60
; 
32'd29480: dataIn1 = 32'd62
; 
32'd29481: dataIn1 = 32'd3
; 
32'd29482: dataIn1 = 32'd4
; 
32'd29483: dataIn1 = 32'd5
; 
32'd29484: dataIn1 = 32'd7
; 
32'd29485: dataIn1 = 32'd9
; 
32'd29486: dataIn1 = 32'd10
; 
32'd29487: dataIn1 = 32'd12
; 
32'd29488: dataIn1 = 32'd18
; 
32'd29489: dataIn1 = 32'd20
; 
32'd29490: dataIn1 = 32'd21
; 
32'd29491: dataIn1 = 32'd23
; 
32'd29492: dataIn1 = 32'd24
; 
32'd29493: dataIn1 = 32'd25
; 
32'd29494: dataIn1 = 32'd27
; 
32'd29495: dataIn1 = 32'd29
; 
32'd29496: dataIn1 = 32'd30
; 
32'd29497: dataIn1 = 32'd31
; 
32'd29498: dataIn1 = 32'd34
; 
32'd29499: dataIn1 = 32'd36
; 
32'd29500: dataIn1 = 32'd39
; 
32'd29501: dataIn1 = 32'd41
; 
32'd29502: dataIn1 = 32'd42
; 
32'd29503: dataIn1 = 32'd43
; 
32'd29504: dataIn1 = 32'd44
; 
32'd29505: dataIn1 = 32'd45
; 
32'd29506: dataIn1 = 32'd48
; 
32'd29507: dataIn1 = 32'd49
; 
32'd29508: dataIn1 = 32'd50
; 
32'd29509: dataIn1 = 32'd53
; 
32'd29510: dataIn1 = 32'd55
; 
32'd29511: dataIn1 = 32'd57
; 
32'd29512: dataIn1 = 32'd63
; 
32'd29513: dataIn1 = 32'd0
; 
32'd29514: dataIn1 = 32'd2
; 
32'd29515: dataIn1 = 32'd4
; 
32'd29516: dataIn1 = 32'd6
; 
32'd29517: dataIn1 = 32'd7
; 
32'd29518: dataIn1 = 32'd8
; 
32'd29519: dataIn1 = 32'd10
; 
32'd29520: dataIn1 = 32'd13
; 
32'd29521: dataIn1 = 32'd14
; 
32'd29522: dataIn1 = 32'd16
; 
32'd29523: dataIn1 = 32'd17
; 
32'd29524: dataIn1 = 32'd18
; 
32'd29525: dataIn1 = 32'd19
; 
32'd29526: dataIn1 = 32'd20
; 
32'd29527: dataIn1 = 32'd23
; 
32'd29528: dataIn1 = 32'd26
; 
32'd29529: dataIn1 = 32'd27
; 
32'd29530: dataIn1 = 32'd30
; 
32'd29531: dataIn1 = 32'd31
; 
32'd29532: dataIn1 = 32'd32
; 
32'd29533: dataIn1 = 32'd36
; 
32'd29534: dataIn1 = 32'd37
; 
32'd29535: dataIn1 = 32'd38
; 
32'd29536: dataIn1 = 32'd40
; 
32'd29537: dataIn1 = 32'd41
; 
32'd29538: dataIn1 = 32'd44
; 
32'd29539: dataIn1 = 32'd46
; 
32'd29540: dataIn1 = 32'd47
; 
32'd29541: dataIn1 = 32'd48
; 
32'd29542: dataIn1 = 32'd49
; 
32'd29543: dataIn1 = 32'd52
; 
32'd29544: dataIn1 = 32'd53
; 
32'd29545: dataIn1 = 32'd54
; 
32'd29546: dataIn1 = 32'd55
; 
32'd29547: dataIn1 = 32'd57
; 
32'd29548: dataIn1 = 32'd58
; 
32'd29549: dataIn1 = 32'd59
; 
32'd29550: dataIn1 = 32'd61
; 
32'd29551: dataIn1 = 32'd0
; 
32'd29552: dataIn1 = 32'd1
; 
32'd29553: dataIn1 = 32'd3
; 
32'd29554: dataIn1 = 32'd4
; 
32'd29555: dataIn1 = 32'd6
; 
32'd29556: dataIn1 = 32'd7
; 
32'd29557: dataIn1 = 32'd8
; 
32'd29558: dataIn1 = 32'd10
; 
32'd29559: dataIn1 = 32'd11
; 
32'd29560: dataIn1 = 32'd12
; 
32'd29561: dataIn1 = 32'd13
; 
32'd29562: dataIn1 = 32'd15
; 
32'd29563: dataIn1 = 32'd16
; 
32'd29564: dataIn1 = 32'd18
; 
32'd29565: dataIn1 = 32'd23
; 
32'd29566: dataIn1 = 32'd26
; 
32'd29567: dataIn1 = 32'd27
; 
32'd29568: dataIn1 = 32'd30
; 
32'd29569: dataIn1 = 32'd31
; 
32'd29570: dataIn1 = 32'd32
; 
32'd29571: dataIn1 = 32'd33
; 
32'd29572: dataIn1 = 32'd34
; 
32'd29573: dataIn1 = 32'd35
; 
32'd29574: dataIn1 = 32'd36
; 
32'd29575: dataIn1 = 32'd37
; 
32'd29576: dataIn1 = 32'd40
; 
32'd29577: dataIn1 = 32'd42
; 
32'd29578: dataIn1 = 32'd44
; 
32'd29579: dataIn1 = 32'd46
; 
32'd29580: dataIn1 = 32'd47
; 
32'd29581: dataIn1 = 32'd48
; 
32'd29582: dataIn1 = 32'd50
; 
32'd29583: dataIn1 = 32'd51
; 
32'd29584: dataIn1 = 32'd53
; 
32'd29585: dataIn1 = 32'd54
; 
32'd29586: dataIn1 = 32'd55
; 
32'd29587: dataIn1 = 32'd57
; 
32'd29588: dataIn1 = 32'd59
; 
32'd29589: dataIn1 = 32'd60
; 
32'd29590: dataIn1 = 32'd61
; 
32'd29591: dataIn1 = 32'd2
; 
32'd29592: dataIn1 = 32'd4
; 
32'd29593: dataIn1 = 32'd6
; 
32'd29594: dataIn1 = 32'd8
; 
32'd29595: dataIn1 = 32'd9
; 
32'd29596: dataIn1 = 32'd10
; 
32'd29597: dataIn1 = 32'd14
; 
32'd29598: dataIn1 = 32'd15
; 
32'd29599: dataIn1 = 32'd16
; 
32'd29600: dataIn1 = 32'd20
; 
32'd29601: dataIn1 = 32'd22
; 
32'd29602: dataIn1 = 32'd23
; 
32'd29603: dataIn1 = 32'd24
; 
32'd29604: dataIn1 = 32'd25
; 
32'd29605: dataIn1 = 32'd27
; 
32'd29606: dataIn1 = 32'd28
; 
32'd29607: dataIn1 = 32'd30
; 
32'd29608: dataIn1 = 32'd32
; 
32'd29609: dataIn1 = 32'd34
; 
32'd29610: dataIn1 = 32'd35
; 
32'd29611: dataIn1 = 32'd41
; 
32'd29612: dataIn1 = 32'd42
; 
32'd29613: dataIn1 = 32'd44
; 
32'd29614: dataIn1 = 32'd45
; 
32'd29615: dataIn1 = 32'd46
; 
32'd29616: dataIn1 = 32'd47
; 
32'd29617: dataIn1 = 32'd48
; 
32'd29618: dataIn1 = 32'd50
; 
32'd29619: dataIn1 = 32'd54
; 
32'd29620: dataIn1 = 32'd55
; 
32'd29621: dataIn1 = 32'd57
; 
32'd29622: dataIn1 = 32'd58
; 
32'd29623: dataIn1 = 32'd60
; 
32'd29624: dataIn1 = 32'd63
; 
32'd29625: dataIn1 = 32'd0
; 
32'd29626: dataIn1 = 32'd2
; 
32'd29627: dataIn1 = 32'd3
; 
32'd29628: dataIn1 = 32'd6
; 
32'd29629: dataIn1 = 32'd7
; 
32'd29630: dataIn1 = 32'd10
; 
32'd29631: dataIn1 = 32'd11
; 
32'd29632: dataIn1 = 32'd12
; 
32'd29633: dataIn1 = 32'd13
; 
32'd29634: dataIn1 = 32'd15
; 
32'd29635: dataIn1 = 32'd17
; 
32'd29636: dataIn1 = 32'd20
; 
32'd29637: dataIn1 = 32'd22
; 
32'd29638: dataIn1 = 32'd24
; 
32'd29639: dataIn1 = 32'd25
; 
32'd29640: dataIn1 = 32'd28
; 
32'd29641: dataIn1 = 32'd31
; 
32'd29642: dataIn1 = 32'd38
; 
32'd29643: dataIn1 = 32'd41
; 
32'd29644: dataIn1 = 32'd42
; 
32'd29645: dataIn1 = 32'd44
; 
32'd29646: dataIn1 = 32'd45
; 
32'd29647: dataIn1 = 32'd47
; 
32'd29648: dataIn1 = 32'd53
; 
32'd29649: dataIn1 = 32'd55
; 
32'd29650: dataIn1 = 32'd56
; 
32'd29651: dataIn1 = 32'd58
; 
32'd29652: dataIn1 = 32'd61
; 
32'd29653: dataIn1 = 32'd62
; 
32'd29654: dataIn1 = 32'd63
; 
32'd29655: dataIn1 = 32'd1
; 
32'd29656: dataIn1 = 32'd10
; 
32'd29657: dataIn1 = 32'd12
; 
32'd29658: dataIn1 = 32'd13
; 
32'd29659: dataIn1 = 32'd14
; 
32'd29660: dataIn1 = 32'd17
; 
32'd29661: dataIn1 = 32'd18
; 
32'd29662: dataIn1 = 32'd19
; 
32'd29663: dataIn1 = 32'd20
; 
32'd29664: dataIn1 = 32'd22
; 
32'd29665: dataIn1 = 32'd24
; 
32'd29666: dataIn1 = 32'd26
; 
32'd29667: dataIn1 = 32'd27
; 
32'd29668: dataIn1 = 32'd28
; 
32'd29669: dataIn1 = 32'd29
; 
32'd29670: dataIn1 = 32'd31
; 
32'd29671: dataIn1 = 32'd32
; 
32'd29672: dataIn1 = 32'd34
; 
32'd29673: dataIn1 = 32'd35
; 
32'd29674: dataIn1 = 32'd38
; 
32'd29675: dataIn1 = 32'd39
; 
32'd29676: dataIn1 = 32'd41
; 
32'd29677: dataIn1 = 32'd43
; 
32'd29678: dataIn1 = 32'd44
; 
32'd29679: dataIn1 = 32'd45
; 
32'd29680: dataIn1 = 32'd46
; 
32'd29681: dataIn1 = 32'd48
; 
32'd29682: dataIn1 = 32'd51
; 
32'd29683: dataIn1 = 32'd52
; 
32'd29684: dataIn1 = 32'd55
; 
32'd29685: dataIn1 = 32'd56
; 
32'd29686: dataIn1 = 32'd57
; 
32'd29687: dataIn1 = 32'd58
; 
32'd29688: dataIn1 = 32'd60
; 
32'd29689: dataIn1 = 32'd61
; 
32'd29690: dataIn1 = 32'd62
; 
32'd29691: dataIn1 = 32'd0
; 
32'd29692: dataIn1 = 32'd1
; 
32'd29693: dataIn1 = 32'd2
; 
32'd29694: dataIn1 = 32'd3
; 
32'd29695: dataIn1 = 32'd6
; 
32'd29696: dataIn1 = 32'd9
; 
32'd29697: dataIn1 = 32'd10
; 
32'd29698: dataIn1 = 32'd12
; 
32'd29699: dataIn1 = 32'd13
; 
32'd29700: dataIn1 = 32'd14
; 
32'd29701: dataIn1 = 32'd16
; 
32'd29702: dataIn1 = 32'd20
; 
32'd29703: dataIn1 = 32'd22
; 
32'd29704: dataIn1 = 32'd23
; 
32'd29705: dataIn1 = 32'd27
; 
32'd29706: dataIn1 = 32'd29
; 
32'd29707: dataIn1 = 32'd33
; 
32'd29708: dataIn1 = 32'd34
; 
32'd29709: dataIn1 = 32'd36
; 
32'd29710: dataIn1 = 32'd37
; 
32'd29711: dataIn1 = 32'd38
; 
32'd29712: dataIn1 = 32'd39
; 
32'd29713: dataIn1 = 32'd40
; 
32'd29714: dataIn1 = 32'd41
; 
32'd29715: dataIn1 = 32'd42
; 
32'd29716: dataIn1 = 32'd45
; 
32'd29717: dataIn1 = 32'd46
; 
32'd29718: dataIn1 = 32'd47
; 
32'd29719: dataIn1 = 32'd51
; 
32'd29720: dataIn1 = 32'd52
; 
32'd29721: dataIn1 = 32'd53
; 
32'd29722: dataIn1 = 32'd55
; 
32'd29723: dataIn1 = 32'd58
; 
32'd29724: dataIn1 = 32'd60
; 
32'd29725: dataIn1 = 32'd61
; 
32'd29726: dataIn1 = 32'd62
; 
32'd29727: dataIn1 = 32'd63
; 
32'd29728: dataIn1 = 32'd0
; 
32'd29729: dataIn1 = 32'd6
; 
32'd29730: dataIn1 = 32'd8
; 
32'd29731: dataIn1 = 32'd10
; 
32'd29732: dataIn1 = 32'd11
; 
32'd29733: dataIn1 = 32'd12
; 
32'd29734: dataIn1 = 32'd14
; 
32'd29735: dataIn1 = 32'd15
; 
32'd29736: dataIn1 = 32'd16
; 
32'd29737: dataIn1 = 32'd18
; 
32'd29738: dataIn1 = 32'd19
; 
32'd29739: dataIn1 = 32'd20
; 
32'd29740: dataIn1 = 32'd22
; 
32'd29741: dataIn1 = 32'd23
; 
32'd29742: dataIn1 = 32'd26
; 
32'd29743: dataIn1 = 32'd27
; 
32'd29744: dataIn1 = 32'd28
; 
32'd29745: dataIn1 = 32'd30
; 
32'd29746: dataIn1 = 32'd34
; 
32'd29747: dataIn1 = 32'd35
; 
32'd29748: dataIn1 = 32'd36
; 
32'd29749: dataIn1 = 32'd37
; 
32'd29750: dataIn1 = 32'd38
; 
32'd29751: dataIn1 = 32'd40
; 
32'd29752: dataIn1 = 32'd42
; 
32'd29753: dataIn1 = 32'd46
; 
32'd29754: dataIn1 = 32'd48
; 
32'd29755: dataIn1 = 32'd51
; 
32'd29756: dataIn1 = 32'd52
; 
32'd29757: dataIn1 = 32'd53
; 
32'd29758: dataIn1 = 32'd55
; 
32'd29759: dataIn1 = 32'd56
; 
32'd29760: dataIn1 = 32'd57
; 
32'd29761: dataIn1 = 32'd60
; 
32'd29762: dataIn1 = 32'd63
; 
32'd29763: dataIn1 = 32'd0
; 
32'd29764: dataIn1 = 32'd2
; 
32'd29765: dataIn1 = 32'd3
; 
32'd29766: dataIn1 = 32'd6
; 
32'd29767: dataIn1 = 32'd7
; 
32'd29768: dataIn1 = 32'd10
; 
32'd29769: dataIn1 = 32'd12
; 
32'd29770: dataIn1 = 32'd13
; 
32'd29771: dataIn1 = 32'd15
; 
32'd29772: dataIn1 = 32'd19
; 
32'd29773: dataIn1 = 32'd20
; 
32'd29774: dataIn1 = 32'd21
; 
32'd29775: dataIn1 = 32'd23
; 
32'd29776: dataIn1 = 32'd24
; 
32'd29777: dataIn1 = 32'd25
; 
32'd29778: dataIn1 = 32'd28
; 
32'd29779: dataIn1 = 32'd29
; 
32'd29780: dataIn1 = 32'd30
; 
32'd29781: dataIn1 = 32'd32
; 
32'd29782: dataIn1 = 32'd34
; 
32'd29783: dataIn1 = 32'd35
; 
32'd29784: dataIn1 = 32'd38
; 
32'd29785: dataIn1 = 32'd40
; 
32'd29786: dataIn1 = 32'd44
; 
32'd29787: dataIn1 = 32'd45
; 
32'd29788: dataIn1 = 32'd50
; 
32'd29789: dataIn1 = 32'd51
; 
32'd29790: dataIn1 = 32'd53
; 
32'd29791: dataIn1 = 32'd54
; 
32'd29792: dataIn1 = 32'd58
; 
32'd29793: dataIn1 = 32'd59
; 
32'd29794: dataIn1 = 32'd60
; 
32'd29795: dataIn1 = 32'd63
; 
32'd29796: dataIn1 = 32'd0
; 
32'd29797: dataIn1 = 32'd1
; 
32'd29798: dataIn1 = 32'd2
; 
32'd29799: dataIn1 = 32'd3
; 
32'd29800: dataIn1 = 32'd5
; 
32'd29801: dataIn1 = 32'd9
; 
32'd29802: dataIn1 = 32'd10
; 
32'd29803: dataIn1 = 32'd12
; 
32'd29804: dataIn1 = 32'd18
; 
32'd29805: dataIn1 = 32'd19
; 
32'd29806: dataIn1 = 32'd20
; 
32'd29807: dataIn1 = 32'd23
; 
32'd29808: dataIn1 = 32'd25
; 
32'd29809: dataIn1 = 32'd27
; 
32'd29810: dataIn1 = 32'd30
; 
32'd29811: dataIn1 = 32'd33
; 
32'd29812: dataIn1 = 32'd34
; 
32'd29813: dataIn1 = 32'd35
; 
32'd29814: dataIn1 = 32'd39
; 
32'd29815: dataIn1 = 32'd41
; 
32'd29816: dataIn1 = 32'd44
; 
32'd29817: dataIn1 = 32'd48
; 
32'd29818: dataIn1 = 32'd49
; 
32'd29819: dataIn1 = 32'd52
; 
32'd29820: dataIn1 = 32'd53
; 
32'd29821: dataIn1 = 32'd56
; 
32'd29822: dataIn1 = 32'd58
; 
32'd29823: dataIn1 = 32'd62
; 
32'd29824: dataIn1 = 32'd63
; 
32'd29825: dataIn1 = 32'd0
; 
32'd29826: dataIn1 = 32'd5
; 
32'd29827: dataIn1 = 32'd6
; 
32'd29828: dataIn1 = 32'd10
; 
32'd29829: dataIn1 = 32'd11
; 
32'd29830: dataIn1 = 32'd13
; 
32'd29831: dataIn1 = 32'd14
; 
32'd29832: dataIn1 = 32'd15
; 
32'd29833: dataIn1 = 32'd19
; 
32'd29834: dataIn1 = 32'd20
; 
32'd29835: dataIn1 = 32'd21
; 
32'd29836: dataIn1 = 32'd22
; 
32'd29837: dataIn1 = 32'd23
; 
32'd29838: dataIn1 = 32'd25
; 
32'd29839: dataIn1 = 32'd27
; 
32'd29840: dataIn1 = 32'd28
; 
32'd29841: dataIn1 = 32'd30
; 
32'd29842: dataIn1 = 32'd31
; 
32'd29843: dataIn1 = 32'd36
; 
32'd29844: dataIn1 = 32'd37
; 
32'd29845: dataIn1 = 32'd39
; 
32'd29846: dataIn1 = 32'd40
; 
32'd29847: dataIn1 = 32'd41
; 
32'd29848: dataIn1 = 32'd43
; 
32'd29849: dataIn1 = 32'd44
; 
32'd29850: dataIn1 = 32'd45
; 
32'd29851: dataIn1 = 32'd47
; 
32'd29852: dataIn1 = 32'd51
; 
32'd29853: dataIn1 = 32'd52
; 
32'd29854: dataIn1 = 32'd54
; 
32'd29855: dataIn1 = 32'd55
; 
32'd29856: dataIn1 = 32'd57
; 
32'd29857: dataIn1 = 32'd58
; 
32'd29858: dataIn1 = 32'd63
; 
32'd29859: dataIn1 = 32'd1
; 
32'd29860: dataIn1 = 32'd2
; 
32'd29861: dataIn1 = 32'd3
; 
32'd29862: dataIn1 = 32'd4
; 
32'd29863: dataIn1 = 32'd5
; 
32'd29864: dataIn1 = 32'd7
; 
32'd29865: dataIn1 = 32'd9
; 
32'd29866: dataIn1 = 32'd12
; 
32'd29867: dataIn1 = 32'd15
; 
32'd29868: dataIn1 = 32'd18
; 
32'd29869: dataIn1 = 32'd19
; 
32'd29870: dataIn1 = 32'd20
; 
32'd29871: dataIn1 = 32'd22
; 
32'd29872: dataIn1 = 32'd24
; 
32'd29873: dataIn1 = 32'd25
; 
32'd29874: dataIn1 = 32'd26
; 
32'd29875: dataIn1 = 32'd27
; 
32'd29876: dataIn1 = 32'd29
; 
32'd29877: dataIn1 = 32'd30
; 
32'd29878: dataIn1 = 32'd32
; 
32'd29879: dataIn1 = 32'd34
; 
32'd29880: dataIn1 = 32'd35
; 
32'd29881: dataIn1 = 32'd37
; 
32'd29882: dataIn1 = 32'd39
; 
32'd29883: dataIn1 = 32'd41
; 
32'd29884: dataIn1 = 32'd43
; 
32'd29885: dataIn1 = 32'd44
; 
32'd29886: dataIn1 = 32'd45
; 
32'd29887: dataIn1 = 32'd47
; 
32'd29888: dataIn1 = 32'd48
; 
32'd29889: dataIn1 = 32'd52
; 
32'd29890: dataIn1 = 32'd53
; 
32'd29891: dataIn1 = 32'd54
; 
32'd29892: dataIn1 = 32'd57
; 
32'd29893: dataIn1 = 32'd60
; 
32'd29894: dataIn1 = 32'd62
; 
32'd29895: dataIn1 = 32'd63
; 
32'd29896: dataIn1 = 32'd0
; 
32'd29897: dataIn1 = 32'd1
; 
32'd29898: dataIn1 = 32'd2
; 
32'd29899: dataIn1 = 32'd3
; 
32'd29900: dataIn1 = 32'd4
; 
32'd29901: dataIn1 = 32'd5
; 
32'd29902: dataIn1 = 32'd6
; 
32'd29903: dataIn1 = 32'd7
; 
32'd29904: dataIn1 = 32'd9
; 
32'd29905: dataIn1 = 32'd10
; 
32'd29906: dataIn1 = 32'd11
; 
32'd29907: dataIn1 = 32'd12
; 
32'd29908: dataIn1 = 32'd13
; 
32'd29909: dataIn1 = 32'd16
; 
32'd29910: dataIn1 = 32'd19
; 
32'd29911: dataIn1 = 32'd20
; 
32'd29912: dataIn1 = 32'd23
; 
32'd29913: dataIn1 = 32'd25
; 
32'd29914: dataIn1 = 32'd26
; 
32'd29915: dataIn1 = 32'd27
; 
32'd29916: dataIn1 = 32'd30
; 
32'd29917: dataIn1 = 32'd31
; 
32'd29918: dataIn1 = 32'd36
; 
32'd29919: dataIn1 = 32'd37
; 
32'd29920: dataIn1 = 32'd38
; 
32'd29921: dataIn1 = 32'd39
; 
32'd29922: dataIn1 = 32'd40
; 
32'd29923: dataIn1 = 32'd41
; 
32'd29924: dataIn1 = 32'd42
; 
32'd29925: dataIn1 = 32'd43
; 
32'd29926: dataIn1 = 32'd46
; 
32'd29927: dataIn1 = 32'd47
; 
32'd29928: dataIn1 = 32'd48
; 
32'd29929: dataIn1 = 32'd50
; 
32'd29930: dataIn1 = 32'd54
; 
32'd29931: dataIn1 = 32'd55
; 
32'd29932: dataIn1 = 32'd56
; 
32'd29933: dataIn1 = 32'd57
; 
32'd29934: dataIn1 = 32'd59
; 
32'd29935: dataIn1 = 32'd61
; 
32'd29936: dataIn1 = 32'd62
; 
32'd29937: dataIn1 = 32'd63
; 
32'd29938: dataIn1 = 32'd0
; 
32'd29939: dataIn1 = 32'd2
; 
32'd29940: dataIn1 = 32'd4
; 
32'd29941: dataIn1 = 32'd5
; 
32'd29942: dataIn1 = 32'd6
; 
32'd29943: dataIn1 = 32'd7
; 
32'd29944: dataIn1 = 32'd9
; 
32'd29945: dataIn1 = 32'd10
; 
32'd29946: dataIn1 = 32'd12
; 
32'd29947: dataIn1 = 32'd14
; 
32'd29948: dataIn1 = 32'd17
; 
32'd29949: dataIn1 = 32'd20
; 
32'd29950: dataIn1 = 32'd21
; 
32'd29951: dataIn1 = 32'd22
; 
32'd29952: dataIn1 = 32'd23
; 
32'd29953: dataIn1 = 32'd25
; 
32'd29954: dataIn1 = 32'd27
; 
32'd29955: dataIn1 = 32'd29
; 
32'd29956: dataIn1 = 32'd30
; 
32'd29957: dataIn1 = 32'd31
; 
32'd29958: dataIn1 = 32'd33
; 
32'd29959: dataIn1 = 32'd35
; 
32'd29960: dataIn1 = 32'd39
; 
32'd29961: dataIn1 = 32'd41
; 
32'd29962: dataIn1 = 32'd42
; 
32'd29963: dataIn1 = 32'd43
; 
32'd29964: dataIn1 = 32'd44
; 
32'd29965: dataIn1 = 32'd45
; 
32'd29966: dataIn1 = 32'd46
; 
32'd29967: dataIn1 = 32'd48
; 
32'd29968: dataIn1 = 32'd49
; 
32'd29969: dataIn1 = 32'd51
; 
32'd29970: dataIn1 = 32'd53
; 
32'd29971: dataIn1 = 32'd55
; 
32'd29972: dataIn1 = 32'd56
; 
32'd29973: dataIn1 = 32'd58
; 
32'd29974: dataIn1 = 32'd59
; 
32'd29975: dataIn1 = 32'd60
; 
32'd29976: dataIn1 = 32'd61
; 
32'd29977: dataIn1 = 32'd62
; 
32'd29978: dataIn1 = 32'd63
; 
32'd29979: dataIn1 = 32'd0
; 
32'd29980: dataIn1 = 32'd2
; 
32'd29981: dataIn1 = 32'd3
; 
32'd29982: dataIn1 = 32'd5
; 
32'd29983: dataIn1 = 32'd6
; 
32'd29984: dataIn1 = 32'd7
; 
32'd29985: dataIn1 = 32'd8
; 
32'd29986: dataIn1 = 32'd10
; 
32'd29987: dataIn1 = 32'd11
; 
32'd29988: dataIn1 = 32'd12
; 
32'd29989: dataIn1 = 32'd13
; 
32'd29990: dataIn1 = 32'd16
; 
32'd29991: dataIn1 = 32'd17
; 
32'd29992: dataIn1 = 32'd18
; 
32'd29993: dataIn1 = 32'd20
; 
32'd29994: dataIn1 = 32'd21
; 
32'd29995: dataIn1 = 32'd22
; 
32'd29996: dataIn1 = 32'd26
; 
32'd29997: dataIn1 = 32'd27
; 
32'd29998: dataIn1 = 32'd30
; 
32'd29999: dataIn1 = 32'd33
; 
32'd30000: dataIn1 = 32'd35
; 
32'd30001: dataIn1 = 32'd36
; 
32'd30002: dataIn1 = 32'd37
; 
32'd30003: dataIn1 = 32'd39
; 
32'd30004: dataIn1 = 32'd40
; 
32'd30005: dataIn1 = 32'd42
; 
32'd30006: dataIn1 = 32'd43
; 
32'd30007: dataIn1 = 32'd44
; 
32'd30008: dataIn1 = 32'd45
; 
32'd30009: dataIn1 = 32'd47
; 
32'd30010: dataIn1 = 32'd48
; 
32'd30011: dataIn1 = 32'd49
; 
32'd30012: dataIn1 = 32'd55
; 
32'd30013: dataIn1 = 32'd56
; 
32'd30014: dataIn1 = 32'd61
; 
32'd30015: dataIn1 = 32'd62
; 
32'd30016: dataIn1 = 32'd1
; 
32'd30017: dataIn1 = 32'd5
; 
32'd30018: dataIn1 = 32'd6
; 
32'd30019: dataIn1 = 32'd8
; 
32'd30020: dataIn1 = 32'd10
; 
32'd30021: dataIn1 = 32'd12
; 
32'd30022: dataIn1 = 32'd13
; 
32'd30023: dataIn1 = 32'd19
; 
32'd30024: dataIn1 = 32'd20
; 
32'd30025: dataIn1 = 32'd25
; 
32'd30026: dataIn1 = 32'd26
; 
32'd30027: dataIn1 = 32'd28
; 
32'd30028: dataIn1 = 32'd29
; 
32'd30029: dataIn1 = 32'd30
; 
32'd30030: dataIn1 = 32'd31
; 
32'd30031: dataIn1 = 32'd34
; 
32'd30032: dataIn1 = 32'd35
; 
32'd30033: dataIn1 = 32'd36
; 
32'd30034: dataIn1 = 32'd37
; 
32'd30035: dataIn1 = 32'd38
; 
32'd30036: dataIn1 = 32'd39
; 
32'd30037: dataIn1 = 32'd41
; 
32'd30038: dataIn1 = 32'd42
; 
32'd30039: dataIn1 = 32'd44
; 
32'd30040: dataIn1 = 32'd46
; 
32'd30041: dataIn1 = 32'd51
; 
32'd30042: dataIn1 = 32'd54
; 
32'd30043: dataIn1 = 32'd55
; 
32'd30044: dataIn1 = 32'd57
; 
32'd30045: dataIn1 = 32'd58
; 
32'd30046: dataIn1 = 32'd59
; 
32'd30047: dataIn1 = 32'd60
; 
32'd30048: dataIn1 = 32'd63
; 
32'd30049: dataIn1 = 32'd0
; 
32'd30050: dataIn1 = 32'd2
; 
32'd30051: dataIn1 = 32'd4
; 
32'd30052: dataIn1 = 32'd5
; 
32'd30053: dataIn1 = 32'd7
; 
32'd30054: dataIn1 = 32'd8
; 
32'd30055: dataIn1 = 32'd9
; 
32'd30056: dataIn1 = 32'd10
; 
32'd30057: dataIn1 = 32'd12
; 
32'd30058: dataIn1 = 32'd13
; 
32'd30059: dataIn1 = 32'd15
; 
32'd30060: dataIn1 = 32'd18
; 
32'd30061: dataIn1 = 32'd19
; 
32'd30062: dataIn1 = 32'd21
; 
32'd30063: dataIn1 = 32'd25
; 
32'd30064: dataIn1 = 32'd26
; 
32'd30065: dataIn1 = 32'd27
; 
32'd30066: dataIn1 = 32'd28
; 
32'd30067: dataIn1 = 32'd29
; 
32'd30068: dataIn1 = 32'd33
; 
32'd30069: dataIn1 = 32'd34
; 
32'd30070: dataIn1 = 32'd36
; 
32'd30071: dataIn1 = 32'd37
; 
32'd30072: dataIn1 = 32'd38
; 
32'd30073: dataIn1 = 32'd41
; 
32'd30074: dataIn1 = 32'd43
; 
32'd30075: dataIn1 = 32'd45
; 
32'd30076: dataIn1 = 32'd46
; 
32'd30077: dataIn1 = 32'd48
; 
32'd30078: dataIn1 = 32'd49
; 
32'd30079: dataIn1 = 32'd52
; 
32'd30080: dataIn1 = 32'd54
; 
32'd30081: dataIn1 = 32'd55
; 
32'd30082: dataIn1 = 32'd56
; 
32'd30083: dataIn1 = 32'd57
; 
32'd30084: dataIn1 = 32'd62
; 
32'd30085: dataIn1 = 32'd63
; 
32'd30086: dataIn1 = 32'd0
; 
32'd30087: dataIn1 = 32'd2
; 
32'd30088: dataIn1 = 32'd3
; 
32'd30089: dataIn1 = 32'd4
; 
32'd30090: dataIn1 = 32'd8
; 
32'd30091: dataIn1 = 32'd9
; 
32'd30092: dataIn1 = 32'd11
; 
32'd30093: dataIn1 = 32'd12
; 
32'd30094: dataIn1 = 32'd14
; 
32'd30095: dataIn1 = 32'd15
; 
32'd30096: dataIn1 = 32'd16
; 
32'd30097: dataIn1 = 32'd17
; 
32'd30098: dataIn1 = 32'd20
; 
32'd30099: dataIn1 = 32'd21
; 
32'd30100: dataIn1 = 32'd23
; 
32'd30101: dataIn1 = 32'd25
; 
32'd30102: dataIn1 = 32'd27
; 
32'd30103: dataIn1 = 32'd28
; 
32'd30104: dataIn1 = 32'd30
; 
32'd30105: dataIn1 = 32'd34
; 
32'd30106: dataIn1 = 32'd36
; 
32'd30107: dataIn1 = 32'd37
; 
32'd30108: dataIn1 = 32'd39
; 
32'd30109: dataIn1 = 32'd40
; 
32'd30110: dataIn1 = 32'd41
; 
32'd30111: dataIn1 = 32'd43
; 
32'd30112: dataIn1 = 32'd44
; 
32'd30113: dataIn1 = 32'd48
; 
32'd30114: dataIn1 = 32'd49
; 
32'd30115: dataIn1 = 32'd50
; 
32'd30116: dataIn1 = 32'd52
; 
32'd30117: dataIn1 = 32'd54
; 
32'd30118: dataIn1 = 32'd56
; 
32'd30119: dataIn1 = 32'd58
; 
32'd30120: dataIn1 = 32'd61
; 
32'd30121: dataIn1 = 32'd62
; 
32'd30122: dataIn1 = 32'd0
; 
32'd30123: dataIn1 = 32'd1
; 
32'd30124: dataIn1 = 32'd2
; 
32'd30125: dataIn1 = 32'd4
; 
32'd30126: dataIn1 = 32'd5
; 
32'd30127: dataIn1 = 32'd6
; 
32'd30128: dataIn1 = 32'd7
; 
32'd30129: dataIn1 = 32'd8
; 
32'd30130: dataIn1 = 32'd10
; 
32'd30131: dataIn1 = 32'd11
; 
32'd30132: dataIn1 = 32'd12
; 
32'd30133: dataIn1 = 32'd14
; 
32'd30134: dataIn1 = 32'd15
; 
32'd30135: dataIn1 = 32'd16
; 
32'd30136: dataIn1 = 32'd19
; 
32'd30137: dataIn1 = 32'd21
; 
32'd30138: dataIn1 = 32'd22
; 
32'd30139: dataIn1 = 32'd24
; 
32'd30140: dataIn1 = 32'd25
; 
32'd30141: dataIn1 = 32'd28
; 
32'd30142: dataIn1 = 32'd30
; 
32'd30143: dataIn1 = 32'd31
; 
32'd30144: dataIn1 = 32'd33
; 
32'd30145: dataIn1 = 32'd36
; 
32'd30146: dataIn1 = 32'd38
; 
32'd30147: dataIn1 = 32'd39
; 
32'd30148: dataIn1 = 32'd44
; 
32'd30149: dataIn1 = 32'd45
; 
32'd30150: dataIn1 = 32'd46
; 
32'd30151: dataIn1 = 32'd47
; 
32'd30152: dataIn1 = 32'd48
; 
32'd30153: dataIn1 = 32'd51
; 
32'd30154: dataIn1 = 32'd52
; 
32'd30155: dataIn1 = 32'd54
; 
32'd30156: dataIn1 = 32'd58
; 
32'd30157: dataIn1 = 32'd60
; 
32'd30158: dataIn1 = 32'd61
; 
32'd30159: dataIn1 = 32'd1
; 
32'd30160: dataIn1 = 32'd2
; 
32'd30161: dataIn1 = 32'd4
; 
32'd30162: dataIn1 = 32'd5
; 
32'd30163: dataIn1 = 32'd6
; 
32'd30164: dataIn1 = 32'd7
; 
32'd30165: dataIn1 = 32'd9
; 
32'd30166: dataIn1 = 32'd11
; 
32'd30167: dataIn1 = 32'd13
; 
32'd30168: dataIn1 = 32'd14
; 
32'd30169: dataIn1 = 32'd15
; 
32'd30170: dataIn1 = 32'd17
; 
32'd30171: dataIn1 = 32'd18
; 
32'd30172: dataIn1 = 32'd19
; 
32'd30173: dataIn1 = 32'd20
; 
32'd30174: dataIn1 = 32'd21
; 
32'd30175: dataIn1 = 32'd26
; 
32'd30176: dataIn1 = 32'd28
; 
32'd30177: dataIn1 = 32'd29
; 
32'd30178: dataIn1 = 32'd30
; 
32'd30179: dataIn1 = 32'd31
; 
32'd30180: dataIn1 = 32'd36
; 
32'd30181: dataIn1 = 32'd38
; 
32'd30182: dataIn1 = 32'd41
; 
32'd30183: dataIn1 = 32'd44
; 
32'd30184: dataIn1 = 32'd46
; 
32'd30185: dataIn1 = 32'd51
; 
32'd30186: dataIn1 = 32'd52
; 
32'd30187: dataIn1 = 32'd54
; 
32'd30188: dataIn1 = 32'd55
; 
32'd30189: dataIn1 = 32'd57
; 
32'd30190: dataIn1 = 32'd58
; 
32'd30191: dataIn1 = 32'd59
; 
32'd30192: dataIn1 = 32'd0
; 
32'd30193: dataIn1 = 32'd1
; 
32'd30194: dataIn1 = 32'd5
; 
32'd30195: dataIn1 = 32'd6
; 
32'd30196: dataIn1 = 32'd7
; 
32'd30197: dataIn1 = 32'd11
; 
32'd30198: dataIn1 = 32'd12
; 
32'd30199: dataIn1 = 32'd15
; 
32'd30200: dataIn1 = 32'd16
; 
32'd30201: dataIn1 = 32'd17
; 
32'd30202: dataIn1 = 32'd18
; 
32'd30203: dataIn1 = 32'd19
; 
32'd30204: dataIn1 = 32'd21
; 
32'd30205: dataIn1 = 32'd24
; 
32'd30206: dataIn1 = 32'd25
; 
32'd30207: dataIn1 = 32'd26
; 
32'd30208: dataIn1 = 32'd28
; 
32'd30209: dataIn1 = 32'd30
; 
32'd30210: dataIn1 = 32'd31
; 
32'd30211: dataIn1 = 32'd32
; 
32'd30212: dataIn1 = 32'd34
; 
32'd30213: dataIn1 = 32'd37
; 
32'd30214: dataIn1 = 32'd40
; 
32'd30215: dataIn1 = 32'd42
; 
32'd30216: dataIn1 = 32'd43
; 
32'd30217: dataIn1 = 32'd44
; 
32'd30218: dataIn1 = 32'd49
; 
32'd30219: dataIn1 = 32'd50
; 
32'd30220: dataIn1 = 32'd51
; 
32'd30221: dataIn1 = 32'd52
; 
32'd30222: dataIn1 = 32'd54
; 
32'd30223: dataIn1 = 32'd55
; 
32'd30224: dataIn1 = 32'd57
; 
32'd30225: dataIn1 = 32'd58
; 
32'd30226: dataIn1 = 32'd62
; 
32'd30227: dataIn1 = 32'd63
; 
32'd30228: dataIn1 = 32'd; 
32'd30229: dataIn1 = 32'd; 
32'd30230: dataIn1 = 32'd; 
32'd30231: dataIn1 = 32'd; 
32'd30232: dataIn1 = 32'd; 
32'd30233: dataIn1 = 32'd; 
32'd30234: dataIn1 = 32'd; 
32'd30235: dataIn1 = 32'd; 
32'd30236: dataIn1 = 32'd; 
32'd30237: dataIn1 = 32'd; 
32'd30238: dataIn1 = 32'd; 
32'd30239: dataIn1 = 32'd; 
32'd30240: dataIn1 = 32'd; 
32'd30241: dataIn1 = 32'd; 
32'd30242: dataIn1 = 32'd; 
32'd30243: dataIn1 = 32'd; 
32'd30244: dataIn1 = 32'd; 
32'd30245: dataIn1 = 32'd; 
32'd30246: dataIn1 = 32'd; 
32'd30247: dataIn1 = 32'd; 
32'd30248: dataIn1 = 32'd; 
32'd30249: dataIn1 = 32'd; 
32'd30250: dataIn1 = 32'd; 
32'd30251: dataIn1 = 32'd; 
32'd30252: dataIn1 = 32'd; 
32'd30253: dataIn1 = 32'd; 
32'd30254: dataIn1 = 32'd; 
32'd30255: dataIn1 = 32'd; 
32'd30256: dataIn1 = 32'd; 
32'd30257: dataIn1 = 32'd; 
32'd30258: dataIn1 = 32'd; 
32'd30259: dataIn1 = 32'd; 
32'd30260: dataIn1 = 32'd; 
32'd30261: dataIn1 = 32'd; 
32'd30262: dataIn1 = 32'd; 
32'd30263: dataIn1 = 32'd; 
32'd30264: dataIn1 = 32'd; 
32'd30265: dataIn1 = 32'd; 
32'd30266: dataIn1 = 32'd; 
32'd30267: dataIn1 = 32'd; 
32'd30268: dataIn1 = 32'd; 
32'd30269: dataIn1 = 32'd; 
32'd30270: dataIn1 = 32'd; 
32'd30271: dataIn1 = 32'd; 
32'd30272: dataIn1 = 32'd; 
32'd30273: dataIn1 = 32'd; 
32'd30274: dataIn1 = 32'd; 
32'd30275: dataIn1 = 32'd; 
32'd30276: dataIn1 = 32'd; 
32'd30277: dataIn1 = 32'd; 
32'd30278: dataIn1 = 32'd; 
32'd30279: dataIn1 = 32'd; 
32'd30280: dataIn1 = 32'd; 
32'd30281: dataIn1 = 32'd; 
32'd30282: dataIn1 = 32'd; 
32'd30283: dataIn1 = 32'd; 
32'd30284: dataIn1 = 32'd; 
32'd30285: dataIn1 = 32'd; 
32'd30286: dataIn1 = 32'd; 
32'd30287: dataIn1 = 32'd; 
32'd30288: dataIn1 = 32'd; 
32'd30289: dataIn1 = 32'd; 
32'd30290: dataIn1 = 32'd; 
32'd30291: dataIn1 = 32'd; 
32'd30292: dataIn1 = 32'd; 
32'd30293: dataIn1 = 32'd; 
32'd30294: dataIn1 = 32'd; 
32'd30295: dataIn1 = 32'd; 
32'd30296: dataIn1 = 32'd; 
32'd30297: dataIn1 = 32'd; 
32'd30298: dataIn1 = 32'd; 
32'd30299: dataIn1 = 32'd; 
32'd30300: dataIn1 = 32'd; 
32'd30301: dataIn1 = 32'd; 
32'd30302: dataIn1 = 32'd; 
32'd30303: dataIn1 = 32'd; 
32'd30304: dataIn1 = 32'd; 
32'd30305: dataIn1 = 32'd; 
32'd30306: dataIn1 = 32'd; 
32'd30307: dataIn1 = 32'd; 
32'd30308: dataIn1 = 32'd; 
32'd30309: dataIn1 = 32'd; 
32'd30310: dataIn1 = 32'd; 
32'd30311: dataIn1 = 32'd; 
32'd30312: dataIn1 = 32'd; 
32'd30313: dataIn1 = 32'd; 
32'd30314: dataIn1 = 32'd; 
32'd30315: dataIn1 = 32'd; 
32'd30316: dataIn1 = 32'd; 
32'd30317: dataIn1 = 32'd; 
32'd30318: dataIn1 = 32'd; 
32'd30319: dataIn1 = 32'd; 
32'd30320: dataIn1 = 32'd; 
32'd30321: dataIn1 = 32'd; 
32'd30322: dataIn1 = 32'd; 
32'd30323: dataIn1 = 32'd; 
32'd30324: dataIn1 = 32'd; 
32'd30325: dataIn1 = 32'd; 
32'd30326: dataIn1 = 32'd; 
32'd30327: dataIn1 = 32'd; 
32'd30328: dataIn1 = 32'd; 
32'd30329: dataIn1 = 32'd; 
32'd30330: dataIn1 = 32'd; 
32'd30331: dataIn1 = 32'd; 
32'd30332: dataIn1 = 32'd; 
32'd30333: dataIn1 = 32'd; 
32'd30334: dataIn1 = 32'd; 
32'd30335: dataIn1 = 32'd; 
32'd30336: dataIn1 = 32'd; 
32'd30337: dataIn1 = 32'd; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd29; 
32'd3: dataIn2 = 32'd55; 
32'd4: dataIn2 = 32'd10; 
32'd5: dataIn2 = 32'd63; 
32'd6: dataIn2 = 32'd23; 
32'd7: dataIn2 = 32'd80; 
32'd8: dataIn2 = 32'd20; 
32'd9: dataIn2 = 32'd39; 
32'd10: dataIn2 = 32'd7; 
32'd11: dataIn2 = 32'd4; 
32'd12: dataIn2 = 32'd82; 
32'd13: dataIn2 = 32'd61; 
32'd14: dataIn2 = 32'd22; 
32'd15: dataIn2 = 32'd14; 
32'd16: dataIn2 = 32'd76; 
32'd17: dataIn2 = 32'd46; 
32'd18: dataIn2 = 32'd75; 
32'd19: dataIn2 = 32'd74; 
32'd20: dataIn2 = 32'd7; 
32'd21: dataIn2 = 32'd65; 
32'd22: dataIn2 = 32'd58; 
32'd23: dataIn2 = 32'd62; 
32'd24: dataIn2 = 32'd100; 
32'd25: dataIn2 = 32'd22; 
32'd26: dataIn2 = 32'd28; 
32'd27: dataIn2 = 32'd62; 
32'd28: dataIn2 = 32'd10; 
32'd29: dataIn2 = 32'd12; 
32'd30: dataIn2 = 32'd46; 
32'd31: dataIn2 = 32'd83; 
32'd32: dataIn2 = 32'd29; 
32'd33: dataIn2 = 32'd1; 
32'd34: dataIn2 = 32'd50; 
32'd35: dataIn2 = 32'd33; 
32'd36: dataIn2 = 32'd18; 
32'd37: dataIn2 = 32'd71; 
32'd38: dataIn2 = 32'd88; 
32'd39: dataIn2 = 32'd4; 
32'd40: dataIn2 = 32'd11; 
32'd41: dataIn2 = 32'd93; 
32'd42: dataIn2 = 32'd76; 
32'd43: dataIn2 = 32'd42; 
32'd44: dataIn2 = 32'd12; 
32'd45: dataIn2 = 32'd25; 
32'd46: dataIn2 = 32'd12; 
32'd47: dataIn2 = 32'd52; 
32'd48: dataIn2 = 32'd38; 
32'd49: dataIn2 = 32'd80; 
32'd50: dataIn2 = 32'd1; 
32'd51: dataIn2 = 32'd28; 
32'd52: dataIn2 = 32'd3; 
32'd53: dataIn2 = 32'd75; 
32'd54: dataIn2 = 32'd62; 
32'd55: dataIn2 = 32'd18; 
32'd56: dataIn2 = 32'd5; 
32'd57: dataIn2 = 32'd10; 
32'd58: dataIn2 = 32'd39; 
32'd59: dataIn2 = 32'd59; 
32'd60: dataIn2 = 32'd96; 
32'd61: dataIn2 = 32'd57; 
32'd62: dataIn2 = 32'd45; 
32'd63: dataIn2 = 32'd6; 
32'd64: dataIn2 = 32'd90; 
32'd65: dataIn2 = 32'd74; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd330: dataIn2 = 32'd80; 
32'd331: dataIn2 = 32'd68; 
32'd332: dataIn2 = 32'd28; 
32'd333: dataIn2 = 32'd60; 
32'd334: dataIn2 = 32'd27; 
32'd335: dataIn2 = 32'd11; 
32'd336: dataIn2 = 32'd0; 
32'd337: dataIn2 = 32'd65; 
32'd338: dataIn2 = 32'd5; 
32'd339: dataIn2 = 32'd15; 
32'd340: dataIn2 = 32'd55; 
32'd341: dataIn2 = 32'd6; 
32'd342: dataIn2 = 32'd25; 
32'd343: dataIn2 = 32'd61; 
32'd344: dataIn2 = 32'd4; 
32'd345: dataIn2 = 32'd83; 
32'd346: dataIn2 = 32'd94; 
32'd347: dataIn2 = 32'd47; 
32'd348: dataIn2 = 32'd24; 
32'd349: dataIn2 = 32'd88; 
32'd350: dataIn2 = 32'd25; 
32'd351: dataIn2 = 32'd23; 
32'd352: dataIn2 = 32'd73; 
32'd353: dataIn2 = 32'd12; 
32'd354: dataIn2 = 32'd81; 
32'd355: dataIn2 = 32'd83; 
32'd356: dataIn2 = 32'd23; 
32'd357: dataIn2 = 32'd91; 
32'd358: dataIn2 = 32'd91; 
32'd359: dataIn2 = 32'd38; 
32'd360: dataIn2 = 32'd40; 
32'd361: dataIn2 = 32'd58; 
32'd362: dataIn2 = 32'd11; 
32'd363: dataIn2 = 32'd83; 
32'd364: dataIn2 = 32'd13; 
32'd365: dataIn2 = 32'd48; 
32'd366: dataIn2 = 32'd49; 
32'd367: dataIn2 = 32'd56; 
32'd368: dataIn2 = 32'd86; 
32'd369: dataIn2 = 32'd61; 
32'd370: dataIn2 = 32'd40; 
32'd371: dataIn2 = 32'd18; 
32'd372: dataIn2 = 32'd27; 
32'd373: dataIn2 = 32'd63; 
32'd374: dataIn2 = 32'd79; 
32'd375: dataIn2 = 32'd50; 
32'd376: dataIn2 = 32'd11; 
32'd377: dataIn2 = 32'd74; 
32'd378: dataIn2 = 32'd81; 
32'd379: dataIn2 = 32'd65; 
32'd380: dataIn2 = 32'd6; 
32'd381: dataIn2 = 32'd69; 
32'd382: dataIn2 = 32'd8; 
32'd383: dataIn2 = 32'd14; 
32'd384: dataIn2 = 32'd39; 
32'd385: dataIn2 = 32'd22; 
32'd386: dataIn2 = 32'd84; 
32'd387: dataIn2 = 32'd51; 
32'd388: dataIn2 = 32'd78; 
32'd389: dataIn2 = 32'd38; 
32'd390: dataIn2 = 32'd73; 
32'd391: dataIn2 = 32'd35; 
32'd392: dataIn2 = 32'd68; 
32'd393: dataIn2 = 32'd52; 
32'd394: dataIn2 = 32'd91; 
32'd395: dataIn2 = 32'd70; 
32'd396: dataIn2 = 32'd11; 
32'd397: dataIn2 = 32'd26; 
32'd398: dataIn2 = 32'd42; 
32'd399: dataIn2 = 32'd44; 
32'd400: dataIn2 = 32'd83; 
32'd401: dataIn2 = 32'd16; 
32'd402: dataIn2 = 32'd93; 
32'd403: dataIn2 = 32'd74; 
32'd404: dataIn2 = 32'd99; 
32'd405: dataIn2 = 32'd93; 
32'd406: dataIn2 = 32'd41; 
32'd407: dataIn2 = 32'd9; 
32'd408: dataIn2 = 32'd14; 
32'd409: dataIn2 = 32'd25; 
32'd410: dataIn2 = 32'd43; 
32'd411: dataIn2 = 32'd26; 
32'd412: dataIn2 = 32'd2; 
32'd413: dataIn2 = 32'd0; 
32'd414: dataIn2 = 32'd2; 
32'd415: dataIn2 = 32'd82; 
32'd416: dataIn2 = 32'd33; 
32'd417: dataIn2 = 32'd80; 
32'd418: dataIn2 = 32'd90; 
32'd419: dataIn2 = 32'd69; 
32'd420: dataIn2 = 32'd52; 
32'd421: dataIn2 = 32'd80; 
32'd422: dataIn2 = 32'd60; 
32'd423: dataIn2 = 32'd38; 
32'd424: dataIn2 = 32'd51; 
32'd425: dataIn2 = 32'd95; 
32'd426: dataIn2 = 32'd58; 
32'd427: dataIn2 = 32'd29; 
32'd428: dataIn2 = 32'd81; 
32'd429: dataIn2 = 32'd23; 
32'd430: dataIn2 = 32'd81; 
32'd431: dataIn2 = 32'd71; 
32'd432: dataIn2 = 32'd5; 
32'd433: dataIn2 = 32'd64; 
32'd434: dataIn2 = 32'd20; 
32'd435: dataIn2 = 32'd86; 
32'd436: dataIn2 = 32'd85; 
32'd437: dataIn2 = 32'd36; 
32'd438: dataIn2 = 32'd24; 
32'd439: dataIn2 = 32'd54; 
32'd440: dataIn2 = 32'd75; 
32'd441: dataIn2 = 32'd69; 
32'd442: dataIn2 = 32'd36; 
32'd443: dataIn2 = 32'd13; 
32'd444: dataIn2 = 32'd63; 
32'd445: dataIn2 = 32'd80; 
32'd446: dataIn2 = 32'd85; 
32'd447: dataIn2 = 32'd89; 
32'd448: dataIn2 = 32'd56; 
32'd449: dataIn2 = 32'd89; 
32'd450: dataIn2 = 32'd48; 
32'd451: dataIn2 = 32'd22; 
32'd452: dataIn2 = 32'd55; 
32'd453: dataIn2 = 32'd72; 
32'd454: dataIn2 = 32'd55; 
32'd455: dataIn2 = 32'd79; 
32'd456: dataIn2 = 32'd80; 
32'd457: dataIn2 = 32'd2; 
32'd458: dataIn2 = 32'd26; 
32'd459: dataIn2 = 32'd48; 
32'd460: dataIn2 = 32'd30; 
32'd461: dataIn2 = 32'd71; 
32'd462: dataIn2 = 32'd91; 
32'd463: dataIn2 = 32'd63; 
32'd464: dataIn2 = 32'd45; 
32'd465: dataIn2 = 32'd64; 
32'd466: dataIn2 = 32'd21; 
32'd467: dataIn2 = 32'd90; 
32'd468: dataIn2 = 32'd0; 
32'd469: dataIn2 = 32'd40; 
32'd470: dataIn2 = 32'd94; 
32'd471: dataIn2 = 32'd53; 
32'd472: dataIn2 = 32'd52; 
32'd473: dataIn2 = 32'd51; 
32'd474: dataIn2 = 32'd54; 
32'd475: dataIn2 = 32'd73; 
32'd476: dataIn2 = 32'd91; 
32'd477: dataIn2 = 32'd99; 
32'd478: dataIn2 = 32'd44; 
32'd479: dataIn2 = 32'd44; 
32'd480: dataIn2 = 32'd16; 
32'd481: dataIn2 = 32'd1; 
32'd482: dataIn2 = 32'd55; 
32'd483: dataIn2 = 32'd38; 
32'd484: dataIn2 = 32'd21; 
32'd485: dataIn2 = 32'd90; 
32'd486: dataIn2 = 32'd27; 
32'd487: dataIn2 = 32'd76; 
32'd488: dataIn2 = 32'd8; 
32'd489: dataIn2 = 32'd84; 
32'd490: dataIn2 = 32'd36; 
32'd491: dataIn2 = 32'd24; 
32'd492: dataIn2 = 32'd64; 
32'd493: dataIn2 = 32'd75; 
32'd494: dataIn2 = 32'd71; 
32'd495: dataIn2 = 32'd87; 
32'd496: dataIn2 = 32'd72; 
32'd497: dataIn2 = 32'd51; 
32'd498: dataIn2 = 32'd97; 
32'd499: dataIn2 = 32'd15; 
32'd500: dataIn2 = 32'd33; 
32'd501: dataIn2 = 32'd50; 
32'd502: dataIn2 = 32'd10; 
32'd503: dataIn2 = 32'd68; 
32'd504: dataIn2 = 32'd36; 
32'd505: dataIn2 = 32'd1; 
32'd506: dataIn2 = 32'd60; 
32'd507: dataIn2 = 32'd67; 
32'd508: dataIn2 = 32'd16; 
32'd509: dataIn2 = 32'd74; 
32'd510: dataIn2 = 32'd5; 
32'd511: dataIn2 = 32'd63; 
32'd512: dataIn2 = 32'd80; 
32'd513: dataIn2 = 32'd24; 
32'd514: dataIn2 = 32'd9; 
32'd515: dataIn2 = 32'd57; 
32'd516: dataIn2 = 32'd8; 
32'd517: dataIn2 = 32'd47; 
32'd518: dataIn2 = 32'd43; 
32'd519: dataIn2 = 32'd95; 
32'd520: dataIn2 = 32'd51; 
32'd521: dataIn2 = 32'd25; 
32'd522: dataIn2 = 32'd40; 
32'd523: dataIn2 = 32'd2; 
32'd524: dataIn2 = 32'd1; 
32'd525: dataIn2 = 32'd21; 
32'd526: dataIn2 = 32'd97; 
32'd527: dataIn2 = 32'd8; 
32'd528: dataIn2 = 32'd10; 
32'd529: dataIn2 = 32'd72; 
32'd530: dataIn2 = 32'd9; 
32'd531: dataIn2 = 32'd43; 
32'd532: dataIn2 = 32'd78; 
32'd533: dataIn2 = 32'd97; 
32'd534: dataIn2 = 32'd32; 
32'd535: dataIn2 = 32'd17; 
32'd536: dataIn2 = 32'd78; 
32'd537: dataIn2 = 32'd33; 
32'd538: dataIn2 = 32'd61; 
32'd539: dataIn2 = 32'd79; 
32'd540: dataIn2 = 32'd62; 
32'd541: dataIn2 = 32'd14; 
32'd542: dataIn2 = 32'd17; 
32'd543: dataIn2 = 32'd88; 
32'd544: dataIn2 = 32'd75; 
32'd545: dataIn2 = 32'd73; 
32'd546: dataIn2 = 32'd1; 
32'd547: dataIn2 = 32'd54; 
32'd548: dataIn2 = 32'd67; 
32'd549: dataIn2 = 32'd27; 
32'd550: dataIn2 = 32'd71; 
32'd551: dataIn2 = 32'd8; 
32'd552: dataIn2 = 32'd34; 
32'd553: dataIn2 = 32'd32; 
32'd554: dataIn2 = 32'd55; 
32'd555: dataIn2 = 32'd80; 
32'd556: dataIn2 = 32'd38; 
32'd557: dataIn2 = 32'd10; 
32'd558: dataIn2 = 32'd26; 
32'd559: dataIn2 = 32'd93; 
32'd560: dataIn2 = 32'd43; 
32'd561: dataIn2 = 32'd43; 
32'd562: dataIn2 = 32'd66; 
32'd563: dataIn2 = 32'd41; 
32'd564: dataIn2 = 32'd68; 
32'd565: dataIn2 = 32'd16; 
32'd566: dataIn2 = 32'd77; 
32'd567: dataIn2 = 32'd83; 
32'd568: dataIn2 = 32'd11; 
32'd569: dataIn2 = 32'd5; 
32'd570: dataIn2 = 32'd35; 
32'd571: dataIn2 = 32'd23; 
32'd572: dataIn2 = 32'd78; 
32'd573: dataIn2 = 32'd81; 
32'd574: dataIn2 = 32'd76; 
32'd575: dataIn2 = 32'd97; 
32'd576: dataIn2 = 32'd26; 
32'd577: dataIn2 = 32'd18; 
32'd578: dataIn2 = 32'd65; 
32'd579: dataIn2 = 32'd85; 
32'd580: dataIn2 = 32'd29; 
32'd581: dataIn2 = 32'd0; 
32'd582: dataIn2 = 32'd74; 
32'd583: dataIn2 = 32'd18; 
32'd584: dataIn2 = 32'd62; 
32'd585: dataIn2 = 32'd92; 
32'd586: dataIn2 = 32'd96; 
32'd587: dataIn2 = 32'd47; 
32'd588: dataIn2 = 32'd69; 
32'd589: dataIn2 = 32'd93; 
32'd590: dataIn2 = 32'd31; 
32'd591: dataIn2 = 32'd66; 
32'd592: dataIn2 = 32'd20; 
32'd593: dataIn2 = 32'd53; 
32'd594: dataIn2 = 32'd29; 
32'd595: dataIn2 = 32'd26; 
32'd596: dataIn2 = 32'd84; 
32'd597: dataIn2 = 32'd67; 
32'd598: dataIn2 = 32'd20; 
32'd599: dataIn2 = 32'd76; 
32'd600: dataIn2 = 32'd64; 
32'd601: dataIn2 = 32'd16; 
32'd602: dataIn2 = 32'd2; 
32'd603: dataIn2 = 32'd96; 
32'd604: dataIn2 = 32'd97; 
32'd605: dataIn2 = 32'd39; 
32'd606: dataIn2 = 32'd36; 
32'd607: dataIn2 = 32'd97; 
32'd608: dataIn2 = 32'd99; 
32'd609: dataIn2 = 32'd69; 
32'd610: dataIn2 = 32'd17; 
32'd611: dataIn2 = 32'd90; 
32'd612: dataIn2 = 32'd36; 
32'd613: dataIn2 = 32'd7; 
32'd614: dataIn2 = 32'd75; 
32'd615: dataIn2 = 32'd4; 
32'd616: dataIn2 = 32'd69; 
32'd617: dataIn2 = 32'd6; 
32'd618: dataIn2 = 32'd23; 
32'd619: dataIn2 = 32'd24; 
32'd620: dataIn2 = 32'd5; 
32'd621: dataIn2 = 32'd58; 
32'd622: dataIn2 = 32'd57; 
32'd623: dataIn2 = 32'd92; 
32'd624: dataIn2 = 32'd50; 
32'd625: dataIn2 = 32'd43; 
32'd626: dataIn2 = 32'd50; 
32'd627: dataIn2 = 32'd92; 
32'd628: dataIn2 = 32'd17; 
32'd629: dataIn2 = 32'd50; 
32'd630: dataIn2 = 32'd34; 
32'd631: dataIn2 = 32'd81; 
32'd632: dataIn2 = 32'd28; 
32'd633: dataIn2 = 32'd72; 
32'd634: dataIn2 = 32'd18; 
32'd635: dataIn2 = 32'd5; 
32'd636: dataIn2 = 32'd61; 
32'd637: dataIn2 = 32'd0; 
32'd638: dataIn2 = 32'd100; 
32'd639: dataIn2 = 32'd83; 
32'd640: dataIn2 = 32'd26; 
32'd641: dataIn2 = 32'd74; 
32'd642: dataIn2 = 32'd16; 
32'd643: dataIn2 = 32'd31; 
32'd644: dataIn2 = 32'd87; 
32'd645: dataIn2 = 32'd95; 
32'd646: dataIn2 = 32'd64; 
32'd647: dataIn2 = 32'd80; 
32'd648: dataIn2 = 32'd82; 
32'd649: dataIn2 = 32'd89; 
32'd650: dataIn2 = 32'd89; 
32'd651: dataIn2 = 32'd68; 
32'd652: dataIn2 = 32'd68; 
32'd653: dataIn2 = 32'd59; 
32'd654: dataIn2 = 32'd17; 
32'd655: dataIn2 = 32'd70; 
32'd656: dataIn2 = 32'd18; 
32'd657: dataIn2 = 32'd22; 
32'd658: dataIn2 = 32'd29; 
32'd659: dataIn2 = 32'd32; 
32'd660: dataIn2 = 32'd73; 
32'd661: dataIn2 = 32'd55; 
32'd662: dataIn2 = 32'd93; 
32'd663: dataIn2 = 32'd48; 
32'd664: dataIn2 = 32'd43; 
32'd665: dataIn2 = 32'd97; 
32'd666: dataIn2 = 32'd32; 
32'd667: dataIn2 = 32'd87; 
32'd668: dataIn2 = 32'd40; 
32'd669: dataIn2 = 32'd98; 
32'd670: dataIn2 = 32'd30; 
32'd671: dataIn2 = 32'd99; 
32'd672: dataIn2 = 32'd51; 
32'd673: dataIn2 = 32'd82; 
32'd674: dataIn2 = 32'd47; 
32'd675: dataIn2 = 32'd76; 
32'd676: dataIn2 = 32'd51; 
32'd677: dataIn2 = 32'd53; 
32'd678: dataIn2 = 32'd22; 
32'd679: dataIn2 = 32'd44; 
32'd680: dataIn2 = 32'd83; 
32'd681: dataIn2 = 32'd95; 
32'd682: dataIn2 = 32'd7; 
32'd683: dataIn2 = 32'd37; 
32'd684: dataIn2 = 32'd9; 
32'd685: dataIn2 = 32'd35; 
32'd686: dataIn2 = 32'd56; 
32'd687: dataIn2 = 32'd2; 
32'd688: dataIn2 = 32'd8; 
32'd689: dataIn2 = 32'd4; 
32'd690: dataIn2 = 32'd74; 
32'd691: dataIn2 = 32'd78; 
32'd692: dataIn2 = 32'd39; 
32'd693: dataIn2 = 32'd99; 
32'd694: dataIn2 = 32'd39; 
32'd695: dataIn2 = 32'd9; 
32'd696: dataIn2 = 32'd47; 
32'd697: dataIn2 = 32'd23; 
32'd698: dataIn2 = 32'd2; 
32'd699: dataIn2 = 32'd68; 
32'd700: dataIn2 = 32'd71; 
32'd701: dataIn2 = 32'd50; 
32'd702: dataIn2 = 32'd54; 
32'd703: dataIn2 = 32'd65; 
32'd704: dataIn2 = 32'd9; 
32'd705: dataIn2 = 32'd97; 
32'd706: dataIn2 = 32'd60; 
32'd707: dataIn2 = 32'd56; 
32'd708: dataIn2 = 32'd82; 
32'd709: dataIn2 = 32'd92; 
32'd710: dataIn2 = 32'd95; 
32'd711: dataIn2 = 32'd95; 
32'd712: dataIn2 = 32'd38; 
32'd713: dataIn2 = 32'd48; 
32'd714: dataIn2 = 32'd59; 
32'd715: dataIn2 = 32'd95; 
32'd716: dataIn2 = 32'd57; 
32'd717: dataIn2 = 32'd99; 
32'd718: dataIn2 = 32'd40; 
32'd719: dataIn2 = 32'd67; 
32'd720: dataIn2 = 32'd76; 
32'd721: dataIn2 = 32'd99; 
32'd722: dataIn2 = 32'd86; 
32'd723: dataIn2 = 32'd41; 
32'd724: dataIn2 = 32'd15; 
32'd725: dataIn2 = 32'd12; 
32'd726: dataIn2 = 32'd74; 
32'd727: dataIn2 = 32'd94; 
32'd728: dataIn2 = 32'd93; 
32'd729: dataIn2 = 32'd76; 
32'd730: dataIn2 = 32'd47; 
32'd731: dataIn2 = 32'd49; 
32'd732: dataIn2 = 32'd50; 
32'd733: dataIn2 = 32'd41; 
32'd734: dataIn2 = 32'd60; 
32'd735: dataIn2 = 32'd62; 
32'd736: dataIn2 = 32'd81; 
32'd737: dataIn2 = 32'd15; 
32'd738: dataIn2 = 32'd71; 
32'd739: dataIn2 = 32'd5; 
32'd740: dataIn2 = 32'd47; 
32'd741: dataIn2 = 32'd29; 
32'd742: dataIn2 = 32'd55; 
32'd743: dataIn2 = 32'd41; 
32'd744: dataIn2 = 32'd6; 
32'd745: dataIn2 = 32'd47; 
32'd746: dataIn2 = 32'd11; 
32'd747: dataIn2 = 32'd94; 
32'd748: dataIn2 = 32'd3; 
32'd749: dataIn2 = 32'd41; 
32'd750: dataIn2 = 32'd57; 
32'd751: dataIn2 = 32'd60; 
32'd752: dataIn2 = 32'd6; 
32'd753: dataIn2 = 32'd40; 
32'd754: dataIn2 = 32'd30; 
32'd755: dataIn2 = 32'd75; 
32'd756: dataIn2 = 32'd86; 
32'd757: dataIn2 = 32'd91; 
32'd758: dataIn2 = 32'd43; 
32'd759: dataIn2 = 32'd50; 
32'd760: dataIn2 = 32'd52; 
32'd761: dataIn2 = 32'd74; 
32'd762: dataIn2 = 32'd58; 
32'd763: dataIn2 = 32'd42; 
32'd764: dataIn2 = 32'd36; 
32'd765: dataIn2 = 32'd39; 
32'd766: dataIn2 = 32'd82; 
32'd767: dataIn2 = 32'd74; 
32'd768: dataIn2 = 32'd55; 
32'd769: dataIn2 = 32'd53; 
32'd770: dataIn2 = 32'd38; 
32'd771: dataIn2 = 32'd92; 
32'd772: dataIn2 = 32'd60; 
32'd773: dataIn2 = 32'd90; 
32'd774: dataIn2 = 32'd14; 
32'd775: dataIn2 = 32'd69; 
32'd776: dataIn2 = 32'd34; 
32'd777: dataIn2 = 32'd82; 
32'd778: dataIn2 = 32'd1; 
32'd779: dataIn2 = 32'd9; 
32'd780: dataIn2 = 32'd80; 
32'd781: dataIn2 = 32'd20; 
32'd782: dataIn2 = 32'd87; 
32'd783: dataIn2 = 32'd71; 
32'd784: dataIn2 = 32'd87; 
32'd785: dataIn2 = 32'd97; 
32'd786: dataIn2 = 32'd83; 
32'd787: dataIn2 = 32'd51; 
32'd788: dataIn2 = 32'd27; 
32'd789: dataIn2 = 32'd90; 
32'd790: dataIn2 = 32'd61; 
32'd791: dataIn2 = 32'd71; 
32'd792: dataIn2 = 32'd82; 
32'd793: dataIn2 = 32'd3; 
32'd794: dataIn2 = 32'd14; 
32'd795: dataIn2 = 32'd21; 
32'd796: dataIn2 = 32'd49; 
32'd797: dataIn2 = 32'd97; 
32'd798: dataIn2 = 32'd36; 
32'd799: dataIn2 = 32'd21; 
32'd800: dataIn2 = 32'd35; 
32'd801: dataIn2 = 32'd6; 
32'd802: dataIn2 = 32'd55; 
32'd803: dataIn2 = 32'd48; 
32'd804: dataIn2 = 32'd52; 
32'd805: dataIn2 = 32'd93; 
32'd806: dataIn2 = 32'd18; 
32'd807: dataIn2 = 32'd3; 
32'd808: dataIn2 = 32'd16; 
32'd809: dataIn2 = 32'd9; 
32'd810: dataIn2 = 32'd48; 
32'd811: dataIn2 = 32'd81; 
32'd812: dataIn2 = 32'd63; 
32'd813: dataIn2 = 32'd12; 
32'd814: dataIn2 = 32'd9; 
32'd815: dataIn2 = 32'd47; 
32'd816: dataIn2 = 32'd42; 
32'd817: dataIn2 = 32'd26; 
32'd818: dataIn2 = 32'd13; 
32'd819: dataIn2 = 32'd43; 
32'd820: dataIn2 = 32'd65; 
32'd821: dataIn2 = 32'd28; 
32'd822: dataIn2 = 32'd38; 
32'd823: dataIn2 = 32'd79; 
32'd824: dataIn2 = 32'd69; 
32'd825: dataIn2 = 32'd38; 
32'd826: dataIn2 = 32'd94; 
32'd827: dataIn2 = 32'd3; 
32'd828: dataIn2 = 32'd65; 
32'd829: dataIn2 = 32'd85; 
32'd830: dataIn2 = 32'd97; 
32'd831: dataIn2 = 32'd70; 
32'd832: dataIn2 = 32'd16; 
32'd833: dataIn2 = 32'd20; 
32'd834: dataIn2 = 32'd32; 
32'd835: dataIn2 = 32'd74; 
32'd836: dataIn2 = 32'd46; 
32'd837: dataIn2 = 32'd4; 
32'd838: dataIn2 = 32'd65; 
32'd839: dataIn2 = 32'd55; 
32'd840: dataIn2 = 32'd23; 
32'd841: dataIn2 = 32'd87; 
32'd842: dataIn2 = 32'd11; 
32'd843: dataIn2 = 32'd19; 
32'd844: dataIn2 = 32'd10; 
32'd845: dataIn2 = 32'd78; 
32'd846: dataIn2 = 32'd82; 
32'd847: dataIn2 = 32'd90; 
32'd848: dataIn2 = 32'd24; 
32'd849: dataIn2 = 32'd50; 
32'd850: dataIn2 = 32'd32; 
32'd851: dataIn2 = 32'd81; 
32'd852: dataIn2 = 32'd15; 
32'd853: dataIn2 = 32'd26; 
32'd854: dataIn2 = 32'd67; 
32'd855: dataIn2 = 32'd71; 
32'd856: dataIn2 = 32'd32; 
32'd857: dataIn2 = 32'd90; 
32'd858: dataIn2 = 32'd32; 
32'd859: dataIn2 = 32'd47; 
32'd860: dataIn2 = 32'd85; 
32'd861: dataIn2 = 32'd26; 
32'd862: dataIn2 = 32'd5; 
32'd863: dataIn2 = 32'd79; 
32'd864: dataIn2 = 32'd33; 
32'd865: dataIn2 = 32'd49; 
32'd866: dataIn2 = 32'd19; 
32'd867: dataIn2 = 32'd9; 
32'd868: dataIn2 = 32'd99; 
32'd869: dataIn2 = 32'd88; 
32'd870: dataIn2 = 32'd18; 
32'd871: dataIn2 = 32'd25; 
32'd872: dataIn2 = 32'd66; 
32'd873: dataIn2 = 32'd78; 
32'd874: dataIn2 = 32'd79; 
32'd875: dataIn2 = 32'd82; 
32'd876: dataIn2 = 32'd74; 
32'd877: dataIn2 = 32'd75; 
32'd878: dataIn2 = 32'd21; 
32'd879: dataIn2 = 32'd16; 
32'd880: dataIn2 = 32'd90; 
32'd881: dataIn2 = 32'd60; 
32'd882: dataIn2 = 32'd64; 
32'd883: dataIn2 = 32'd94; 
32'd884: dataIn2 = 32'd21; 
32'd885: dataIn2 = 32'd44; 
32'd886: dataIn2 = 32'd34; 
32'd887: dataIn2 = 32'd40; 
32'd888: dataIn2 = 32'd58; 
32'd889: dataIn2 = 32'd53; 
32'd890: dataIn2 = 32'd72; 
32'd891: dataIn2 = 32'd1; 
32'd892: dataIn2 = 32'd75; 
32'd893: dataIn2 = 32'd37; 
32'd894: dataIn2 = 32'd53; 
32'd895: dataIn2 = 32'd53; 
32'd896: dataIn2 = 32'd14; 
32'd897: dataIn2 = 32'd89; 
32'd898: dataIn2 = 32'd23; 
32'd899: dataIn2 = 32'd63; 
32'd900: dataIn2 = 32'd99; 
32'd901: dataIn2 = 32'd43; 
32'd902: dataIn2 = 32'd62; 
32'd903: dataIn2 = 32'd1; 
32'd904: dataIn2 = 32'd79; 
32'd905: dataIn2 = 32'd82; 
32'd906: dataIn2 = 32'd17; 
32'd907: dataIn2 = 32'd29; 
32'd908: dataIn2 = 32'd48; 
32'd909: dataIn2 = 32'd99; 
32'd910: dataIn2 = 32'd16; 
32'd911: dataIn2 = 32'd99; 
32'd912: dataIn2 = 32'd77; 
32'd913: dataIn2 = 32'd6; 
32'd914: dataIn2 = 32'd18; 
32'd915: dataIn2 = 32'd62; 
32'd916: dataIn2 = 32'd63; 
32'd917: dataIn2 = 32'd99; 
32'd918: dataIn2 = 32'd93; 
32'd919: dataIn2 = 32'd62; 
32'd920: dataIn2 = 32'd72; 
32'd921: dataIn2 = 32'd51; 
32'd922: dataIn2 = 32'd7; 
32'd923: dataIn2 = 32'd93; 
32'd924: dataIn2 = 32'd22; 
32'd925: dataIn2 = 32'd91; 
32'd926: dataIn2 = 32'd100; 
32'd927: dataIn2 = 32'd20; 
32'd928: dataIn2 = 32'd24; 
32'd929: dataIn2 = 32'd67; 
32'd930: dataIn2 = 32'd11; 
32'd931: dataIn2 = 32'd25; 
32'd932: dataIn2 = 32'd18; 
32'd933: dataIn2 = 32'd34; 
32'd934: dataIn2 = 32'd45; 
32'd935: dataIn2 = 32'd50; 
32'd936: dataIn2 = 32'd12; 
32'd937: dataIn2 = 32'd86; 
32'd938: dataIn2 = 32'd14; 
32'd939: dataIn2 = 32'd72; 
32'd940: dataIn2 = 32'd83; 
32'd941: dataIn2 = 32'd80; 
32'd942: dataIn2 = 32'd21; 
32'd943: dataIn2 = 32'd34; 
32'd944: dataIn2 = 32'd99; 
32'd945: dataIn2 = 32'd13; 
32'd946: dataIn2 = 32'd85; 
32'd947: dataIn2 = 32'd90; 
32'd948: dataIn2 = 32'd63; 
32'd949: dataIn2 = 32'd30; 
32'd950: dataIn2 = 32'd35; 
32'd951: dataIn2 = 32'd27; 
32'd952: dataIn2 = 32'd63; 
32'd953: dataIn2 = 32'd25; 
32'd954: dataIn2 = 32'd49; 
32'd955: dataIn2 = 32'd58; 
32'd956: dataIn2 = 32'd21; 
32'd957: dataIn2 = 32'd71; 
32'd958: dataIn2 = 32'd85; 
32'd959: dataIn2 = 32'd71; 
32'd960: dataIn2 = 32'd35; 
32'd961: dataIn2 = 32'd46; 
32'd962: dataIn2 = 32'd75; 
32'd963: dataIn2 = 32'd31; 
32'd964: dataIn2 = 32'd68; 
32'd965: dataIn2 = 32'd8; 
32'd966: dataIn2 = 32'd10; 
32'd967: dataIn2 = 32'd6; 
32'd968: dataIn2 = 32'd24; 
32'd969: dataIn2 = 32'd11; 
32'd970: dataIn2 = 32'd79; 
32'd971: dataIn2 = 32'd33; 
32'd972: dataIn2 = 32'd11; 
32'd973: dataIn2 = 32'd31; 
32'd974: dataIn2 = 32'd62; 
32'd975: dataIn2 = 32'd29; 
32'd976: dataIn2 = 32'd9; 
32'd977: dataIn2 = 32'd81; 
32'd978: dataIn2 = 32'd27; 
32'd979: dataIn2 = 32'd29; 
32'd980: dataIn2 = 32'd77; 
32'd981: dataIn2 = 32'd41; 
32'd982: dataIn2 = 32'd17; 
32'd983: dataIn2 = 32'd16; 
32'd984: dataIn2 = 32'd83; 
32'd985: dataIn2 = 32'd33; 
32'd986: dataIn2 = 32'd57; 
32'd987: dataIn2 = 32'd88; 
32'd988: dataIn2 = 32'd37; 
32'd989: dataIn2 = 32'd49; 
32'd990: dataIn2 = 32'd62; 
32'd991: dataIn2 = 32'd86; 
32'd992: dataIn2 = 32'd30; 
32'd993: dataIn2 = 32'd46; 
32'd994: dataIn2 = 32'd54; 
32'd995: dataIn2 = 32'd95; 
32'd996: dataIn2 = 32'd88; 
32'd997: dataIn2 = 32'd69; 
32'd998: dataIn2 = 32'd43; 
32'd999: dataIn2 = 32'd1; 
32'd1000: dataIn2 = 32'd87; 
32'd1001: dataIn2 = 32'd21; 
32'd1002: dataIn2 = 32'd75; 
32'd1003: dataIn2 = 32'd49; 
32'd1004: dataIn2 = 32'd73; 
32'd1005: dataIn2 = 32'd80; 
32'd1006: dataIn2 = 32'd41; 
32'd1007: dataIn2 = 32'd75; 
32'd1008: dataIn2 = 32'd13; 
32'd1009: dataIn2 = 32'd98; 
32'd1010: dataIn2 = 32'd25; 
32'd1011: dataIn2 = 32'd15; 
32'd1012: dataIn2 = 32'd66; 
32'd1013: dataIn2 = 32'd62; 
32'd1014: dataIn2 = 32'd78; 
32'd1015: dataIn2 = 32'd14; 
32'd1016: dataIn2 = 32'd56; 
32'd1017: dataIn2 = 32'd75; 
32'd1018: dataIn2 = 32'd85; 
32'd1019: dataIn2 = 32'd46; 
32'd1020: dataIn2 = 32'd57; 
32'd1021: dataIn2 = 32'd4; 
32'd1022: dataIn2 = 32'd95; 
32'd1023: dataIn2 = 32'd59; 
32'd1024: dataIn2 = 32'd70; 
32'd1025: dataIn2 = 32'd27; 
32'd1026: dataIn2 = 32'd15; 
32'd1027: dataIn2 = 32'd56; 
32'd1028: dataIn2 = 32'd16; 
32'd1029: dataIn2 = 32'd35; 
32'd1030: dataIn2 = 32'd10; 
32'd1031: dataIn2 = 32'd98; 
32'd1032: dataIn2 = 32'd6; 
32'd1033: dataIn2 = 32'd71; 
32'd1034: dataIn2 = 32'd82; 
32'd1035: dataIn2 = 32'd35; 
32'd1036: dataIn2 = 32'd60; 
32'd1037: dataIn2 = 32'd95; 
32'd1038: dataIn2 = 32'd76; 
32'd1039: dataIn2 = 32'd40; 
32'd1040: dataIn2 = 32'd63; 
32'd1041: dataIn2 = 32'd61; 
32'd1042: dataIn2 = 32'd67; 
32'd1043: dataIn2 = 32'd51; 
32'd1044: dataIn2 = 32'd39; 
32'd1045: dataIn2 = 32'd7; 
32'd1046: dataIn2 = 32'd97; 
32'd1047: dataIn2 = 32'd96; 
32'd1048: dataIn2 = 32'd20; 
32'd1049: dataIn2 = 32'd37; 
32'd1050: dataIn2 = 32'd88; 
32'd1051: dataIn2 = 32'd21; 
32'd1052: dataIn2 = 32'd13; 
32'd1053: dataIn2 = 32'd45; 
32'd1054: dataIn2 = 32'd25; 
32'd1055: dataIn2 = 32'd88; 
32'd1056: dataIn2 = 32'd25; 
32'd1057: dataIn2 = 32'd0; 
32'd1058: dataIn2 = 32'd24; 
32'd1059: dataIn2 = 32'd90; 
32'd1060: dataIn2 = 32'd33; 
32'd1061: dataIn2 = 32'd51; 
32'd1062: dataIn2 = 32'd68; 
32'd1063: dataIn2 = 32'd13; 
32'd1064: dataIn2 = 32'd37; 
32'd1065: dataIn2 = 32'd77; 
32'd1066: dataIn2 = 32'd100; 
32'd1067: dataIn2 = 32'd61; 
32'd1068: dataIn2 = 32'd69; 
32'd1069: dataIn2 = 32'd12; 
32'd1070: dataIn2 = 32'd4; 
32'd1071: dataIn2 = 32'd15; 
32'd1072: dataIn2 = 32'd76; 
32'd1073: dataIn2 = 32'd82; 
32'd1074: dataIn2 = 32'd80; 
32'd1075: dataIn2 = 32'd28; 
32'd1076: dataIn2 = 32'd42; 
32'd1077: dataIn2 = 32'd80; 
32'd1078: dataIn2 = 32'd90; 
32'd1079: dataIn2 = 32'd74; 
32'd1080: dataIn2 = 32'd83; 
32'd1081: dataIn2 = 32'd45; 
32'd1082: dataIn2 = 32'd47; 
32'd1083: dataIn2 = 32'd46; 
32'd1084: dataIn2 = 32'd13; 
32'd1085: dataIn2 = 32'd71; 
32'd1086: dataIn2 = 32'd89; 
32'd1087: dataIn2 = 32'd80; 
32'd1088: dataIn2 = 32'd52; 
32'd1089: dataIn2 = 32'd23; 
32'd1090: dataIn2 = 32'd88; 
32'd1091: dataIn2 = 32'd19; 
32'd1092: dataIn2 = 32'd6; 
32'd1093: dataIn2 = 32'd27; 
32'd1094: dataIn2 = 32'd90; 
32'd1095: dataIn2 = 32'd81; 
32'd1096: dataIn2 = 32'd62; 
32'd1097: dataIn2 = 32'd47; 
32'd1098: dataIn2 = 32'd4; 
32'd1099: dataIn2 = 32'd82; 
32'd1100: dataIn2 = 32'd97; 
32'd1101: dataIn2 = 32'd70; 
32'd1102: dataIn2 = 32'd24; 
32'd1103: dataIn2 = 32'd25; 
32'd1104: dataIn2 = 32'd0; 
32'd1105: dataIn2 = 32'd99; 
32'd1106: dataIn2 = 32'd92; 
32'd1107: dataIn2 = 32'd83; 
32'd1108: dataIn2 = 32'd33; 
32'd1109: dataIn2 = 32'd62; 
32'd1110: dataIn2 = 32'd94; 
32'd1111: dataIn2 = 32'd60; 
32'd1112: dataIn2 = 32'd44; 
32'd1113: dataIn2 = 32'd78; 
32'd1114: dataIn2 = 32'd44; 
32'd1115: dataIn2 = 32'd90; 
32'd1116: dataIn2 = 32'd43; 
32'd1117: dataIn2 = 32'd75; 
32'd1118: dataIn2 = 32'd38; 
32'd1119: dataIn2 = 32'd21; 
32'd1120: dataIn2 = 32'd53; 
32'd1121: dataIn2 = 32'd37; 
32'd1122: dataIn2 = 32'd99; 
32'd1123: dataIn2 = 32'd23; 
32'd1124: dataIn2 = 32'd35; 
32'd1125: dataIn2 = 32'd13; 
32'd1126: dataIn2 = 32'd17; 
32'd1127: dataIn2 = 32'd63; 
32'd1128: dataIn2 = 32'd63; 
32'd1129: dataIn2 = 32'd12; 
32'd1130: dataIn2 = 32'd84; 
32'd1131: dataIn2 = 32'd49; 
32'd1132: dataIn2 = 32'd90; 
32'd1133: dataIn2 = 32'd97; 
32'd1134: dataIn2 = 32'd23; 
32'd1135: dataIn2 = 32'd92; 
32'd1136: dataIn2 = 32'd82; 
32'd1137: dataIn2 = 32'd4; 
32'd1138: dataIn2 = 32'd33; 
32'd1139: dataIn2 = 32'd54; 
32'd1140: dataIn2 = 32'd7; 
32'd1141: dataIn2 = 32'd31; 
32'd1142: dataIn2 = 32'd49; 
32'd1143: dataIn2 = 32'd84; 
32'd1144: dataIn2 = 32'd45; 
32'd1145: dataIn2 = 32'd76; 
32'd1146: dataIn2 = 32'd82; 
32'd1147: dataIn2 = 32'd41; 
32'd1148: dataIn2 = 32'd34; 
32'd1149: dataIn2 = 32'd93; 
32'd1150: dataIn2 = 32'd55; 
32'd1151: dataIn2 = 32'd2; 
32'd1152: dataIn2 = 32'd40; 
32'd1153: dataIn2 = 32'd2; 
32'd1154: dataIn2 = 32'd82; 
32'd1155: dataIn2 = 32'd63; 
32'd1156: dataIn2 = 32'd52; 
32'd1157: dataIn2 = 32'd3; 
32'd1158: dataIn2 = 32'd2; 
32'd1159: dataIn2 = 32'd56; 
32'd1160: dataIn2 = 32'd29; 
32'd1161: dataIn2 = 32'd48; 
32'd1162: dataIn2 = 32'd19; 
32'd1163: dataIn2 = 32'd94; 
32'd1164: dataIn2 = 32'd73; 
32'd1165: dataIn2 = 32'd99; 
32'd1166: dataIn2 = 32'd55; 
32'd1167: dataIn2 = 32'd36; 
32'd1168: dataIn2 = 32'd74; 
32'd1169: dataIn2 = 32'd24; 
32'd1170: dataIn2 = 32'd75; 
32'd1171: dataIn2 = 32'd82; 
32'd1172: dataIn2 = 32'd91; 
32'd1173: dataIn2 = 32'd40; 
32'd1174: dataIn2 = 32'd76; 
32'd1175: dataIn2 = 32'd77; 
32'd1176: dataIn2 = 32'd73; 
32'd1177: dataIn2 = 32'd62; 
32'd1178: dataIn2 = 32'd95; 
32'd1179: dataIn2 = 32'd41; 
32'd1180: dataIn2 = 32'd94; 
32'd1181: dataIn2 = 32'd90; 
32'd1182: dataIn2 = 32'd15; 
32'd1183: dataIn2 = 32'd28; 
32'd1184: dataIn2 = 32'd89; 
32'd1185: dataIn2 = 32'd5; 
32'd1186: dataIn2 = 32'd83; 
32'd1187: dataIn2 = 32'd39; 
32'd1188: dataIn2 = 32'd80; 
32'd1189: dataIn2 = 32'd40; 
32'd1190: dataIn2 = 32'd84; 
32'd1191: dataIn2 = 32'd99; 
32'd1192: dataIn2 = 32'd56; 
32'd1193: dataIn2 = 32'd9; 
32'd1194: dataIn2 = 32'd60; 
32'd1195: dataIn2 = 32'd98; 
32'd1196: dataIn2 = 32'd87; 
32'd1197: dataIn2 = 32'd86; 
32'd1198: dataIn2 = 32'd44; 
32'd1199: dataIn2 = 32'd18; 
32'd1200: dataIn2 = 32'd19; 
32'd1201: dataIn2 = 32'd52; 
32'd1202: dataIn2 = 32'd10; 
32'd1203: dataIn2 = 32'd48; 
32'd1204: dataIn2 = 32'd28; 
32'd1205: dataIn2 = 32'd7; 
32'd1206: dataIn2 = 32'd94; 
32'd1207: dataIn2 = 32'd87; 
32'd1208: dataIn2 = 32'd11; 
32'd1209: dataIn2 = 32'd50; 
32'd1210: dataIn2 = 32'd69; 
32'd1211: dataIn2 = 32'd43; 
32'd1212: dataIn2 = 32'd43; 
32'd1213: dataIn2 = 32'd80; 
32'd1214: dataIn2 = 32'd62; 
32'd1215: dataIn2 = 32'd36; 
32'd1216: dataIn2 = 32'd23; 
32'd1217: dataIn2 = 32'd28; 
32'd1218: dataIn2 = 32'd40; 
32'd1219: dataIn2 = 32'd37; 
32'd1220: dataIn2 = 32'd85; 
32'd1221: dataIn2 = 32'd62; 
32'd1222: dataIn2 = 32'd87; 
32'd1223: dataIn2 = 32'd12; 
32'd1224: dataIn2 = 32'd94; 
32'd1225: dataIn2 = 32'd53; 
32'd1226: dataIn2 = 32'd38; 
32'd1227: dataIn2 = 32'd13; 
32'd1228: dataIn2 = 32'd32; 
32'd1229: dataIn2 = 32'd76; 
32'd1230: dataIn2 = 32'd12; 
32'd1231: dataIn2 = 32'd65; 
32'd1232: dataIn2 = 32'd20; 
32'd1233: dataIn2 = 32'd40; 
32'd1234: dataIn2 = 32'd40; 
32'd1235: dataIn2 = 32'd60; 
32'd1236: dataIn2 = 32'd63; 
32'd1237: dataIn2 = 32'd53; 
32'd1238: dataIn2 = 32'd33; 
32'd1239: dataIn2 = 32'd23; 
32'd1240: dataIn2 = 32'd85; 
32'd1241: dataIn2 = 32'd87; 
32'd1242: dataIn2 = 32'd16; 
32'd1243: dataIn2 = 32'd11; 
32'd1244: dataIn2 = 32'd38; 
32'd1245: dataIn2 = 32'd13; 
32'd1246: dataIn2 = 32'd14; 
32'd1247: dataIn2 = 32'd58; 
32'd1248: dataIn2 = 32'd71; 
32'd1249: dataIn2 = 32'd65; 
32'd1250: dataIn2 = 32'd5; 
32'd1251: dataIn2 = 32'd71; 
32'd1252: dataIn2 = 32'd39; 
32'd1253: dataIn2 = 32'd69; 
32'd1254: dataIn2 = 32'd58; 
32'd1255: dataIn2 = 32'd15; 
32'd1256: dataIn2 = 32'd13; 
32'd1257: dataIn2 = 32'd5; 
32'd1258: dataIn2 = 32'd37; 
32'd1259: dataIn2 = 32'd56; 
32'd1260: dataIn2 = 32'd93; 
32'd1261: dataIn2 = 32'd2; 
32'd1262: dataIn2 = 32'd80; 
32'd1263: dataIn2 = 32'd70; 
32'd1264: dataIn2 = 32'd51; 
32'd1265: dataIn2 = 32'd70; 
32'd1266: dataIn2 = 32'd8; 
32'd1267: dataIn2 = 32'd28; 
32'd1268: dataIn2 = 32'd42; 
32'd1269: dataIn2 = 32'd91; 
32'd1270: dataIn2 = 32'd6; 
32'd1271: dataIn2 = 32'd0; 
32'd1272: dataIn2 = 32'd59; 
32'd1273: dataIn2 = 32'd23; 
32'd1274: dataIn2 = 32'd39; 
32'd1275: dataIn2 = 32'd45; 
32'd1276: dataIn2 = 32'd33; 
32'd1277: dataIn2 = 32'd1; 
32'd1278: dataIn2 = 32'd45; 
32'd1279: dataIn2 = 32'd11; 
32'd1280: dataIn2 = 32'd40; 
32'd1281: dataIn2 = 32'd96; 
32'd1282: dataIn2 = 32'd37; 
32'd1283: dataIn2 = 32'd8; 
32'd1284: dataIn2 = 32'd7; 
32'd1285: dataIn2 = 32'd56; 
32'd1286: dataIn2 = 32'd37; 
32'd1287: dataIn2 = 32'd58; 
32'd1288: dataIn2 = 32'd19; 
32'd1289: dataIn2 = 32'd30; 
32'd1290: dataIn2 = 32'd1; 
32'd1291: dataIn2 = 32'd60; 
32'd1292: dataIn2 = 32'd24; 
32'd1293: dataIn2 = 32'd1; 
32'd1294: dataIn2 = 32'd41; 
32'd1295: dataIn2 = 32'd39; 
32'd1296: dataIn2 = 32'd46; 
32'd1297: dataIn2 = 32'd1; 
32'd1298: dataIn2 = 32'd63; 
32'd1299: dataIn2 = 32'd64; 
32'd1300: dataIn2 = 32'd80; 
32'd1301: dataIn2 = 32'd71; 
32'd1302: dataIn2 = 32'd0; 
32'd1303: dataIn2 = 32'd32; 
32'd1304: dataIn2 = 32'd69; 
32'd1305: dataIn2 = 32'd13; 
32'd1306: dataIn2 = 32'd72; 
32'd1307: dataIn2 = 32'd18; 
32'd1308: dataIn2 = 32'd34; 
32'd1309: dataIn2 = 32'd76; 
32'd1310: dataIn2 = 32'd81; 
32'd1311: dataIn2 = 32'd33; 
32'd1312: dataIn2 = 32'd19; 
32'd1313: dataIn2 = 32'd86; 
32'd1314: dataIn2 = 32'd81; 
32'd1315: dataIn2 = 32'd26; 
32'd1316: dataIn2 = 32'd33; 
32'd1317: dataIn2 = 32'd59; 
32'd1318: dataIn2 = 32'd77; 
32'd1319: dataIn2 = 32'd64; 
32'd1320: dataIn2 = 32'd58; 
32'd1321: dataIn2 = 32'd88; 
32'd1322: dataIn2 = 32'd82; 
32'd1323: dataIn2 = 32'd21; 
32'd1324: dataIn2 = 32'd56; 
32'd1325: dataIn2 = 32'd71; 
32'd1326: dataIn2 = 32'd17; 
32'd1327: dataIn2 = 32'd77; 
32'd1328: dataIn2 = 32'd56; 
32'd1329: dataIn2 = 32'd12; 
32'd1330: dataIn2 = 32'd70; 
32'd1331: dataIn2 = 32'd5; 
32'd1332: dataIn2 = 32'd23; 
32'd1333: dataIn2 = 32'd92; 
32'd1334: dataIn2 = 32'd50; 
32'd1335: dataIn2 = 32'd70; 
32'd1336: dataIn2 = 32'd23; 
32'd1337: dataIn2 = 32'd9; 
32'd1338: dataIn2 = 32'd52; 
32'd1339: dataIn2 = 32'd5; 
32'd1340: dataIn2 = 32'd78; 
32'd1341: dataIn2 = 32'd4; 
32'd1342: dataIn2 = 32'd81; 
32'd1343: dataIn2 = 32'd72; 
32'd1344: dataIn2 = 32'd14; 
32'd1345: dataIn2 = 32'd17; 
32'd1346: dataIn2 = 32'd94; 
32'd1347: dataIn2 = 32'd62; 
32'd1348: dataIn2 = 32'd33; 
32'd1349: dataIn2 = 32'd67; 
32'd1350: dataIn2 = 32'd17; 
32'd1351: dataIn2 = 32'd58; 
32'd1352: dataIn2 = 32'd92; 
32'd1353: dataIn2 = 32'd5; 
32'd1354: dataIn2 = 32'd63; 
32'd1355: dataIn2 = 32'd20; 
32'd1356: dataIn2 = 32'd11; 
32'd1357: dataIn2 = 32'd43; 
32'd1358: dataIn2 = 32'd92; 
32'd1359: dataIn2 = 32'd83; 
32'd1360: dataIn2 = 32'd14; 
32'd1361: dataIn2 = 32'd89; 
32'd1362: dataIn2 = 32'd7; 
32'd1363: dataIn2 = 32'd65; 
32'd1364: dataIn2 = 32'd40; 
32'd1365: dataIn2 = 32'd49; 
32'd1366: dataIn2 = 32'd50; 
32'd1367: dataIn2 = 32'd50; 
32'd1368: dataIn2 = 32'd42; 
32'd1369: dataIn2 = 32'd79; 
32'd1370: dataIn2 = 32'd37; 
32'd1371: dataIn2 = 32'd34; 
32'd1372: dataIn2 = 32'd93; 
32'd1373: dataIn2 = 32'd10; 
32'd1374: dataIn2 = 32'd22; 
32'd1375: dataIn2 = 32'd35; 
32'd1376: dataIn2 = 32'd27; 
32'd1377: dataIn2 = 32'd24; 
32'd1378: dataIn2 = 32'd49; 
32'd1379: dataIn2 = 32'd12; 
32'd1380: dataIn2 = 32'd69; 
32'd1381: dataIn2 = 32'd55; 
32'd1382: dataIn2 = 32'd4; 
32'd1383: dataIn2 = 32'd98; 
32'd1384: dataIn2 = 32'd89; 
32'd1385: dataIn2 = 32'd11; 
32'd1386: dataIn2 = 32'd56; 
32'd1387: dataIn2 = 32'd63; 
32'd1388: dataIn2 = 32'd34; 
32'd1389: dataIn2 = 32'd62; 
32'd1390: dataIn2 = 32'd5; 
32'd1391: dataIn2 = 32'd55; 
32'd1392: dataIn2 = 32'd63; 
32'd1393: dataIn2 = 32'd8; 
32'd1394: dataIn2 = 32'd82; 
32'd1395: dataIn2 = 32'd86; 
32'd1396: dataIn2 = 32'd54; 
32'd1397: dataIn2 = 32'd39; 
32'd1398: dataIn2 = 32'd31; 
32'd1399: dataIn2 = 32'd0; 
32'd1400: dataIn2 = 32'd82; 
32'd1401: dataIn2 = 32'd38; 
32'd1402: dataIn2 = 32'd36; 
32'd1403: dataIn2 = 32'd25; 
32'd1404: dataIn2 = 32'd58; 
32'd1405: dataIn2 = 32'd70; 
32'd1406: dataIn2 = 32'd9; 
32'd1407: dataIn2 = 32'd89; 
32'd1408: dataIn2 = 32'd35; 
32'd1409: dataIn2 = 32'd82; 
32'd1410: dataIn2 = 32'd44; 
32'd1411: dataIn2 = 32'd27; 
32'd1412: dataIn2 = 32'd61; 
32'd1413: dataIn2 = 32'd97; 
32'd1414: dataIn2 = 32'd82; 
32'd1415: dataIn2 = 32'd10; 
32'd1416: dataIn2 = 32'd89; 
32'd1417: dataIn2 = 32'd95; 
32'd1418: dataIn2 = 32'd22; 
32'd1419: dataIn2 = 32'd34; 
32'd1420: dataIn2 = 32'd20; 
32'd1421: dataIn2 = 32'd0; 
32'd1422: dataIn2 = 32'd89; 
32'd1423: dataIn2 = 32'd28; 
32'd1424: dataIn2 = 32'd46; 
32'd1425: dataIn2 = 32'd43; 
32'd1426: dataIn2 = 32'd23; 
32'd1427: dataIn2 = 32'd23; 
32'd1428: dataIn2 = 32'd61; 
32'd1429: dataIn2 = 32'd70; 
32'd1430: dataIn2 = 32'd48; 
32'd1431: dataIn2 = 32'd74; 
32'd1432: dataIn2 = 32'd51; 
32'd1433: dataIn2 = 32'd61; 
32'd1434: dataIn2 = 32'd96; 
32'd1435: dataIn2 = 32'd46; 
32'd1436: dataIn2 = 32'd28; 
32'd1437: dataIn2 = 32'd25; 
32'd1438: dataIn2 = 32'd19; 
32'd1439: dataIn2 = 32'd95; 
32'd1440: dataIn2 = 32'd68; 
32'd1441: dataIn2 = 32'd55; 
32'd1442: dataIn2 = 32'd77; 
32'd1443: dataIn2 = 32'd59; 
32'd1444: dataIn2 = 32'd60; 
32'd1445: dataIn2 = 32'd44; 
32'd1446: dataIn2 = 32'd29; 
32'd1447: dataIn2 = 32'd92; 
32'd1448: dataIn2 = 32'd64; 
32'd1449: dataIn2 = 32'd35; 
32'd1450: dataIn2 = 32'd50; 
32'd1451: dataIn2 = 32'd74; 
32'd1452: dataIn2 = 32'd70; 
32'd1453: dataIn2 = 32'd12; 
32'd1454: dataIn2 = 32'd57; 
32'd1455: dataIn2 = 32'd61; 
32'd1456: dataIn2 = 32'd81; 
32'd1457: dataIn2 = 32'd45; 
32'd1458: dataIn2 = 32'd47; 
32'd1459: dataIn2 = 32'd10; 
32'd1460: dataIn2 = 32'd13; 
32'd1461: dataIn2 = 32'd25; 
32'd1462: dataIn2 = 32'd10; 
32'd1463: dataIn2 = 32'd99; 
32'd1464: dataIn2 = 32'd25; 
32'd1465: dataIn2 = 32'd50; 
32'd1466: dataIn2 = 32'd65; 
32'd1467: dataIn2 = 32'd71; 
32'd1468: dataIn2 = 32'd34; 
32'd1469: dataIn2 = 32'd10; 
32'd1470: dataIn2 = 32'd96; 
32'd1471: dataIn2 = 32'd13; 
32'd1472: dataIn2 = 32'd31; 
32'd1473: dataIn2 = 32'd71; 
32'd1474: dataIn2 = 32'd90; 
32'd1475: dataIn2 = 32'd30; 
32'd1476: dataIn2 = 32'd84; 
32'd1477: dataIn2 = 32'd45; 
32'd1478: dataIn2 = 32'd45; 
32'd1479: dataIn2 = 32'd70; 
32'd1480: dataIn2 = 32'd62; 
32'd1481: dataIn2 = 32'd91; 
32'd1482: dataIn2 = 32'd80; 
32'd1483: dataIn2 = 32'd73; 
32'd1484: dataIn2 = 32'd75; 
32'd1485: dataIn2 = 32'd18; 
32'd1486: dataIn2 = 32'd6; 
32'd1487: dataIn2 = 32'd95; 
32'd1488: dataIn2 = 32'd76; 
32'd1489: dataIn2 = 32'd27; 
32'd1490: dataIn2 = 32'd76; 
32'd1491: dataIn2 = 32'd77; 
32'd1492: dataIn2 = 32'd10; 
32'd1493: dataIn2 = 32'd97; 
32'd1494: dataIn2 = 32'd36; 
32'd1495: dataIn2 = 32'd76; 
32'd1496: dataIn2 = 32'd91; 
32'd1497: dataIn2 = 32'd0; 
32'd1498: dataIn2 = 32'd39; 
32'd1499: dataIn2 = 32'd93; 
32'd1500: dataIn2 = 32'd92; 
32'd1501: dataIn2 = 32'd83; 
32'd1502: dataIn2 = 32'd40; 
32'd1503: dataIn2 = 32'd57; 
32'd1504: dataIn2 = 32'd31; 
32'd1505: dataIn2 = 32'd91; 
32'd1506: dataIn2 = 32'd40; 
32'd1507: dataIn2 = 32'd24; 
32'd1508: dataIn2 = 32'd37; 
32'd1509: dataIn2 = 32'd60; 
32'd1510: dataIn2 = 32'd3; 
32'd1511: dataIn2 = 32'd49; 
32'd1512: dataIn2 = 32'd18; 
32'd1513: dataIn2 = 32'd89; 
32'd1514: dataIn2 = 32'd84; 
32'd1515: dataIn2 = 32'd45; 
32'd1516: dataIn2 = 32'd87; 
32'd1517: dataIn2 = 32'd31; 
32'd1518: dataIn2 = 32'd100; 
32'd1519: dataIn2 = 32'd50; 
32'd1520: dataIn2 = 32'd23; 
32'd1521: dataIn2 = 32'd86; 
32'd1522: dataIn2 = 32'd8; 
32'd1523: dataIn2 = 32'd39; 
32'd1524: dataIn2 = 32'd85; 
32'd1525: dataIn2 = 32'd4; 
32'd1526: dataIn2 = 32'd27; 
32'd1527: dataIn2 = 32'd38; 
32'd1528: dataIn2 = 32'd36; 
32'd1529: dataIn2 = 32'd14; 
32'd1530: dataIn2 = 32'd20; 
32'd1531: dataIn2 = 32'd73; 
32'd1532: dataIn2 = 32'd20; 
32'd1533: dataIn2 = 32'd13; 
32'd1534: dataIn2 = 32'd64; 
32'd1535: dataIn2 = 32'd62; 
32'd1536: dataIn2 = 32'd81; 
32'd1537: dataIn2 = 32'd39; 
32'd1538: dataIn2 = 32'd8; 
32'd1539: dataIn2 = 32'd77; 
32'd1540: dataIn2 = 32'd59; 
32'd1541: dataIn2 = 32'd21; 
32'd1542: dataIn2 = 32'd39; 
32'd1543: dataIn2 = 32'd16; 
32'd1544: dataIn2 = 32'd34; 
32'd1545: dataIn2 = 32'd17; 
32'd1546: dataIn2 = 32'd72; 
32'd1547: dataIn2 = 32'd8; 
32'd1548: dataIn2 = 32'd63; 
32'd1549: dataIn2 = 32'd100; 
32'd1550: dataIn2 = 32'd31; 
32'd1551: dataIn2 = 32'd92; 
32'd1552: dataIn2 = 32'd47; 
32'd1553: dataIn2 = 32'd11; 
32'd1554: dataIn2 = 32'd33; 
32'd1555: dataIn2 = 32'd54; 
32'd1556: dataIn2 = 32'd86; 
32'd1557: dataIn2 = 32'd19; 
32'd1558: dataIn2 = 32'd71; 
32'd1559: dataIn2 = 32'd62; 
32'd1560: dataIn2 = 32'd93; 
32'd1561: dataIn2 = 32'd61; 
32'd1562: dataIn2 = 32'd93; 
32'd1563: dataIn2 = 32'd51; 
32'd1564: dataIn2 = 32'd67; 
32'd1565: dataIn2 = 32'd81; 
32'd1566: dataIn2 = 32'd27; 
32'd1567: dataIn2 = 32'd90; 
32'd1568: dataIn2 = 32'd6; 
32'd1569: dataIn2 = 32'd54; 
32'd1570: dataIn2 = 32'd55; 
32'd1571: dataIn2 = 32'd60; 
32'd1572: dataIn2 = 32'd16; 
32'd1573: dataIn2 = 32'd57; 
32'd1574: dataIn2 = 32'd74; 
32'd1575: dataIn2 = 32'd24; 
32'd1576: dataIn2 = 32'd50; 
32'd1577: dataIn2 = 32'd46; 
32'd1578: dataIn2 = 32'd33; 
32'd1579: dataIn2 = 32'd6; 
32'd1580: dataIn2 = 32'd45; 
32'd1581: dataIn2 = 32'd29; 
32'd1582: dataIn2 = 32'd41; 
32'd1583: dataIn2 = 32'd62; 
32'd1584: dataIn2 = 32'd42; 
32'd1585: dataIn2 = 32'd33; 
32'd1586: dataIn2 = 32'd46; 
32'd1587: dataIn2 = 32'd39; 
32'd1588: dataIn2 = 32'd62; 
32'd1589: dataIn2 = 32'd44; 
32'd1590: dataIn2 = 32'd60; 
32'd1591: dataIn2 = 32'd75; 
32'd1592: dataIn2 = 32'd80; 
32'd1593: dataIn2 = 32'd9; 
32'd1594: dataIn2 = 32'd100; 
32'd1595: dataIn2 = 32'd42; 
32'd1596: dataIn2 = 32'd63; 
32'd1597: dataIn2 = 32'd31; 
32'd1598: dataIn2 = 32'd35; 
32'd1599: dataIn2 = 32'd20; 
32'd1600: dataIn2 = 32'd23; 
32'd1601: dataIn2 = 32'd27; 
32'd1602: dataIn2 = 32'd4; 
32'd1603: dataIn2 = 32'd75; 
32'd1604: dataIn2 = 32'd72; 
32'd1605: dataIn2 = 32'd44; 
32'd1606: dataIn2 = 32'd70; 
32'd1607: dataIn2 = 32'd65; 
32'd1608: dataIn2 = 32'd96; 
32'd1609: dataIn2 = 32'd4; 
32'd1610: dataIn2 = 32'd22; 
32'd1611: dataIn2 = 32'd9; 
32'd1612: dataIn2 = 32'd77; 
32'd1613: dataIn2 = 32'd64; 
32'd1614: dataIn2 = 32'd10; 
32'd1615: dataIn2 = 32'd91; 
32'd1616: dataIn2 = 32'd13; 
32'd1617: dataIn2 = 32'd20; 
32'd1618: dataIn2 = 32'd22; 
32'd1619: dataIn2 = 32'd83; 
32'd1620: dataIn2 = 32'd72; 
32'd1621: dataIn2 = 32'd87; 
32'd1622: dataIn2 = 32'd72; 
32'd1623: dataIn2 = 32'd48; 
32'd1624: dataIn2 = 32'd40; 
32'd1625: dataIn2 = 32'd48; 
32'd1626: dataIn2 = 32'd2; 
32'd1627: dataIn2 = 32'd30; 
32'd1628: dataIn2 = 32'd60; 
32'd1629: dataIn2 = 32'd25; 
32'd1630: dataIn2 = 32'd95; 
32'd1631: dataIn2 = 32'd1; 
32'd1632: dataIn2 = 32'd31; 
32'd1633: dataIn2 = 32'd48; 
32'd1634: dataIn2 = 32'd86; 
32'd1635: dataIn2 = 32'd81; 
32'd1636: dataIn2 = 32'd6; 
32'd1637: dataIn2 = 32'd39; 
32'd1638: dataIn2 = 32'd12; 
32'd1639: dataIn2 = 32'd44; 
32'd1640: dataIn2 = 32'd50; 
32'd1641: dataIn2 = 32'd100; 
32'd1642: dataIn2 = 32'd66; 
32'd1643: dataIn2 = 32'd3; 
32'd1644: dataIn2 = 32'd93; 
32'd1645: dataIn2 = 32'd9; 
32'd1646: dataIn2 = 32'd30; 
32'd1647: dataIn2 = 32'd87; 
32'd1648: dataIn2 = 32'd0; 
32'd1649: dataIn2 = 32'd31; 
32'd1650: dataIn2 = 32'd40; 
32'd1651: dataIn2 = 32'd84; 
32'd1652: dataIn2 = 32'd52; 
32'd1653: dataIn2 = 32'd25; 
32'd1654: dataIn2 = 32'd4; 
32'd1655: dataIn2 = 32'd48; 
32'd1656: dataIn2 = 32'd44; 
32'd1657: dataIn2 = 32'd42; 
32'd1658: dataIn2 = 32'd12; 
32'd1659: dataIn2 = 32'd67; 
32'd1660: dataIn2 = 32'd91; 
32'd1661: dataIn2 = 32'd13; 
32'd1662: dataIn2 = 32'd91; 
32'd1663: dataIn2 = 32'd71; 
32'd1664: dataIn2 = 32'd73; 
32'd1665: dataIn2 = 32'd76; 
32'd1666: dataIn2 = 32'd91; 
32'd1667: dataIn2 = 32'd31; 
32'd1668: dataIn2 = 32'd5; 
32'd1669: dataIn2 = 32'd99; 
32'd1670: dataIn2 = 32'd15; 
32'd1671: dataIn2 = 32'd60; 
32'd1672: dataIn2 = 32'd100; 
32'd1673: dataIn2 = 32'd74; 
32'd1674: dataIn2 = 32'd97; 
32'd1675: dataIn2 = 32'd15; 
32'd1676: dataIn2 = 32'd12; 
32'd1677: dataIn2 = 32'd52; 
32'd1678: dataIn2 = 32'd68; 
32'd1679: dataIn2 = 32'd36; 
32'd1680: dataIn2 = 32'd77; 
32'd1681: dataIn2 = 32'd85; 
32'd1682: dataIn2 = 32'd35; 
32'd1683: dataIn2 = 32'd92; 
32'd1684: dataIn2 = 32'd92; 
32'd1685: dataIn2 = 32'd40; 
32'd1686: dataIn2 = 32'd57; 
32'd1687: dataIn2 = 32'd76; 
32'd1688: dataIn2 = 32'd41; 
32'd1689: dataIn2 = 32'd83; 
32'd1690: dataIn2 = 32'd72; 
32'd1691: dataIn2 = 32'd64; 
32'd1692: dataIn2 = 32'd3; 
32'd1693: dataIn2 = 32'd78; 
32'd1694: dataIn2 = 32'd61; 
32'd1695: dataIn2 = 32'd43; 
32'd1696: dataIn2 = 32'd31; 
32'd1697: dataIn2 = 32'd18; 
32'd1698: dataIn2 = 32'd99; 
32'd1699: dataIn2 = 32'd99; 
32'd1700: dataIn2 = 32'd88; 
32'd1701: dataIn2 = 32'd52; 
32'd1702: dataIn2 = 32'd73; 
32'd1703: dataIn2 = 32'd26; 
32'd1704: dataIn2 = 32'd7; 
32'd1705: dataIn2 = 32'd5; 
32'd1706: dataIn2 = 32'd33; 
32'd1707: dataIn2 = 32'd12; 
32'd1708: dataIn2 = 32'd99; 
32'd1709: dataIn2 = 32'd72; 
32'd1710: dataIn2 = 32'd58; 
32'd1711: dataIn2 = 32'd91; 
32'd1712: dataIn2 = 32'd19; 
32'd1713: dataIn2 = 32'd2; 
32'd1714: dataIn2 = 32'd24; 
32'd1715: dataIn2 = 32'd86; 
32'd1716: dataIn2 = 32'd48; 
32'd1717: dataIn2 = 32'd86; 
32'd1718: dataIn2 = 32'd35; 
32'd1719: dataIn2 = 32'd81; 
32'd1720: dataIn2 = 32'd12; 
32'd1721: dataIn2 = 32'd76; 
32'd1722: dataIn2 = 32'd61; 
32'd1723: dataIn2 = 32'd75; 
32'd1724: dataIn2 = 32'd81; 
32'd1725: dataIn2 = 32'd18; 
32'd1726: dataIn2 = 32'd78; 
32'd1727: dataIn2 = 32'd42; 
32'd1728: dataIn2 = 32'd7; 
32'd1729: dataIn2 = 32'd87; 
32'd1730: dataIn2 = 32'd75; 
32'd1731: dataIn2 = 32'd53; 
32'd1732: dataIn2 = 32'd62; 
32'd1733: dataIn2 = 32'd65; 
32'd1734: dataIn2 = 32'd30; 
32'd1735: dataIn2 = 32'd23; 
32'd1736: dataIn2 = 32'd98; 
32'd1737: dataIn2 = 32'd87; 
32'd1738: dataIn2 = 32'd96; 
32'd1739: dataIn2 = 32'd80; 
32'd1740: dataIn2 = 32'd99; 
32'd1741: dataIn2 = 32'd0; 
32'd1742: dataIn2 = 32'd27; 
32'd1743: dataIn2 = 32'd9; 
32'd1744: dataIn2 = 32'd16; 
32'd1745: dataIn2 = 32'd79; 
32'd1746: dataIn2 = 32'd59; 
32'd1747: dataIn2 = 32'd45; 
32'd1748: dataIn2 = 32'd10; 
32'd1749: dataIn2 = 32'd5; 
32'd1750: dataIn2 = 32'd19; 
32'd1751: dataIn2 = 32'd21; 
32'd1752: dataIn2 = 32'd93; 
32'd1753: dataIn2 = 32'd22; 
32'd1754: dataIn2 = 32'd96; 
32'd1755: dataIn2 = 32'd43; 
32'd1756: dataIn2 = 32'd96; 
32'd1757: dataIn2 = 32'd62; 
32'd1758: dataIn2 = 32'd45; 
32'd1759: dataIn2 = 32'd90; 
32'd1760: dataIn2 = 32'd19; 
32'd1761: dataIn2 = 32'd61; 
32'd1762: dataIn2 = 32'd45; 
32'd1763: dataIn2 = 32'd85; 
32'd1764: dataIn2 = 32'd15; 
32'd1765: dataIn2 = 32'd48; 
32'd1766: dataIn2 = 32'd82; 
32'd1767: dataIn2 = 32'd10; 
32'd1768: dataIn2 = 32'd39; 
32'd1769: dataIn2 = 32'd30; 
32'd1770: dataIn2 = 32'd77; 
32'd1771: dataIn2 = 32'd34; 
32'd1772: dataIn2 = 32'd0; 
32'd1773: dataIn2 = 32'd44; 
32'd1774: dataIn2 = 32'd96; 
32'd1775: dataIn2 = 32'd34; 
32'd1776: dataIn2 = 32'd70; 
32'd1777: dataIn2 = 32'd22; 
32'd1778: dataIn2 = 32'd48; 
32'd1779: dataIn2 = 32'd12; 
32'd1780: dataIn2 = 32'd49; 
32'd1781: dataIn2 = 32'd17; 
32'd1782: dataIn2 = 32'd79; 
32'd1783: dataIn2 = 32'd6; 
32'd1784: dataIn2 = 32'd58; 
32'd1785: dataIn2 = 32'd89; 
32'd1786: dataIn2 = 32'd10; 
32'd1787: dataIn2 = 32'd32; 
32'd1788: dataIn2 = 32'd93; 
32'd1789: dataIn2 = 32'd78; 
32'd1790: dataIn2 = 32'd38; 
32'd1791: dataIn2 = 32'd48; 
32'd1792: dataIn2 = 32'd45; 
32'd1793: dataIn2 = 32'd5; 
32'd1794: dataIn2 = 32'd96; 
32'd1795: dataIn2 = 32'd73; 
32'd1796: dataIn2 = 32'd11; 
32'd1797: dataIn2 = 32'd49; 
32'd1798: dataIn2 = 32'd42; 
32'd1799: dataIn2 = 32'd10; 
32'd1800: dataIn2 = 32'd83; 
32'd1801: dataIn2 = 32'd88; 
32'd1802: dataIn2 = 32'd7; 
32'd1803: dataIn2 = 32'd93; 
32'd1804: dataIn2 = 32'd49; 
32'd1805: dataIn2 = 32'd74; 
32'd1806: dataIn2 = 32'd89; 
32'd1807: dataIn2 = 32'd48; 
32'd1808: dataIn2 = 32'd48; 
32'd1809: dataIn2 = 32'd79; 
32'd1810: dataIn2 = 32'd62; 
32'd1811: dataIn2 = 32'd55; 
32'd1812: dataIn2 = 32'd12; 
32'd1813: dataIn2 = 32'd0; 
32'd1814: dataIn2 = 32'd96; 
32'd1815: dataIn2 = 32'd1; 
32'd1816: dataIn2 = 32'd69; 
32'd1817: dataIn2 = 32'd7; 
32'd1818: dataIn2 = 32'd66; 
32'd1819: dataIn2 = 32'd85; 
32'd1820: dataIn2 = 32'd28; 
32'd1821: dataIn2 = 32'd96; 
32'd1822: dataIn2 = 32'd56; 
32'd1823: dataIn2 = 32'd49; 
32'd1824: dataIn2 = 32'd29; 
32'd1825: dataIn2 = 32'd95; 
32'd1826: dataIn2 = 32'd43; 
32'd1827: dataIn2 = 32'd66; 
32'd1828: dataIn2 = 32'd57; 
32'd1829: dataIn2 = 32'd61; 
32'd1830: dataIn2 = 32'd88; 
32'd1831: dataIn2 = 32'd43; 
32'd1832: dataIn2 = 32'd92; 
32'd1833: dataIn2 = 32'd21; 
32'd1834: dataIn2 = 32'd96; 
32'd1835: dataIn2 = 32'd66; 
32'd1836: dataIn2 = 32'd80; 
32'd1837: dataIn2 = 32'd16; 
32'd1838: dataIn2 = 32'd81; 
32'd1839: dataIn2 = 32'd44; 
32'd1840: dataIn2 = 32'd79; 
32'd1841: dataIn2 = 32'd94; 
32'd1842: dataIn2 = 32'd86; 
32'd1843: dataIn2 = 32'd92; 
32'd1844: dataIn2 = 32'd86; 
32'd1845: dataIn2 = 32'd81; 
32'd1846: dataIn2 = 32'd35; 
32'd1847: dataIn2 = 32'd49; 
32'd1848: dataIn2 = 32'd97; 
32'd1849: dataIn2 = 32'd52; 
32'd1850: dataIn2 = 32'd86; 
32'd1851: dataIn2 = 32'd10; 
32'd1852: dataIn2 = 32'd79; 
32'd1853: dataIn2 = 32'd66; 
32'd1854: dataIn2 = 32'd68; 
32'd1855: dataIn2 = 32'd51; 
32'd1856: dataIn2 = 32'd22; 
32'd1857: dataIn2 = 32'd4; 
32'd1858: dataIn2 = 32'd59; 
32'd1859: dataIn2 = 32'd36; 
32'd1860: dataIn2 = 32'd7; 
32'd1861: dataIn2 = 32'd46; 
32'd1862: dataIn2 = 32'd26; 
32'd1863: dataIn2 = 32'd91; 
32'd1864: dataIn2 = 32'd79; 
32'd1865: dataIn2 = 32'd26; 
32'd1866: dataIn2 = 32'd93; 
32'd1867: dataIn2 = 32'd23; 
32'd1868: dataIn2 = 32'd8; 
32'd1869: dataIn2 = 32'd53; 
32'd1870: dataIn2 = 32'd39; 
32'd1871: dataIn2 = 32'd86; 
32'd1872: dataIn2 = 32'd33; 
32'd1873: dataIn2 = 32'd22; 
32'd1874: dataIn2 = 32'd5; 
32'd1875: dataIn2 = 32'd37; 
32'd1876: dataIn2 = 32'd22; 
32'd1877: dataIn2 = 32'd54; 
32'd1878: dataIn2 = 32'd36; 
32'd1879: dataIn2 = 32'd28; 
32'd1880: dataIn2 = 32'd36; 
32'd1881: dataIn2 = 32'd12; 
32'd1882: dataIn2 = 32'd71; 
32'd1883: dataIn2 = 32'd15; 
32'd1884: dataIn2 = 32'd63; 
32'd1885: dataIn2 = 32'd61; 
32'd1886: dataIn2 = 32'd73; 
32'd1887: dataIn2 = 32'd17; 
32'd1888: dataIn2 = 32'd56; 
32'd1889: dataIn2 = 32'd73; 
32'd1890: dataIn2 = 32'd52; 
32'd1891: dataIn2 = 32'd98; 
32'd1892: dataIn2 = 32'd46; 
32'd1893: dataIn2 = 32'd49; 
32'd1894: dataIn2 = 32'd31; 
32'd1895: dataIn2 = 32'd80; 
32'd1896: dataIn2 = 32'd38; 
32'd1897: dataIn2 = 32'd3; 
32'd1898: dataIn2 = 32'd23; 
32'd1899: dataIn2 = 32'd48; 
32'd1900: dataIn2 = 32'd73; 
32'd1901: dataIn2 = 32'd28; 
32'd1902: dataIn2 = 32'd92; 
32'd1903: dataIn2 = 32'd71; 
32'd1904: dataIn2 = 32'd2; 
32'd1905: dataIn2 = 32'd94; 
32'd1906: dataIn2 = 32'd71; 
32'd1907: dataIn2 = 32'd55; 
32'd1908: dataIn2 = 32'd11; 
32'd1909: dataIn2 = 32'd87; 
32'd1910: dataIn2 = 32'd15; 
32'd1911: dataIn2 = 32'd36; 
32'd1912: dataIn2 = 32'd13; 
32'd1913: dataIn2 = 32'd49; 
32'd1914: dataIn2 = 32'd0; 
32'd1915: dataIn2 = 32'd44; 
32'd1916: dataIn2 = 32'd8; 
32'd1917: dataIn2 = 32'd52; 
32'd1918: dataIn2 = 32'd58; 
32'd1919: dataIn2 = 32'd17; 
32'd1920: dataIn2 = 32'd21; 
32'd1921: dataIn2 = 32'd85; 
32'd1922: dataIn2 = 32'd98; 
32'd1923: dataIn2 = 32'd10; 
32'd1924: dataIn2 = 32'd56; 
32'd1925: dataIn2 = 32'd39; 
32'd1926: dataIn2 = 32'd37; 
32'd1927: dataIn2 = 32'd60; 
32'd1928: dataIn2 = 32'd2; 
32'd1929: dataIn2 = 32'd60; 
32'd1930: dataIn2 = 32'd59; 
32'd1931: dataIn2 = 32'd99; 
32'd1932: dataIn2 = 32'd97; 
32'd1933: dataIn2 = 32'd73; 
32'd1934: dataIn2 = 32'd27; 
32'd1935: dataIn2 = 32'd48; 
32'd1936: dataIn2 = 32'd37; 
32'd1937: dataIn2 = 32'd34; 
32'd1938: dataIn2 = 32'd56; 
32'd1939: dataIn2 = 32'd56; 
32'd1940: dataIn2 = 32'd52; 
32'd1941: dataIn2 = 32'd31; 
32'd1942: dataIn2 = 32'd97; 
32'd1943: dataIn2 = 32'd34; 
32'd1944: dataIn2 = 32'd16; 
32'd1945: dataIn2 = 32'd35; 
32'd1946: dataIn2 = 32'd84; 
32'd1947: dataIn2 = 32'd76; 
32'd1948: dataIn2 = 32'd74; 
32'd1949: dataIn2 = 32'd32; 
32'd1950: dataIn2 = 32'd2; 
32'd1951: dataIn2 = 32'd14; 
32'd1952: dataIn2 = 32'd39; 
32'd1953: dataIn2 = 32'd24; 
32'd1954: dataIn2 = 32'd100; 
32'd1955: dataIn2 = 32'd91; 
32'd1956: dataIn2 = 32'd30; 
32'd1957: dataIn2 = 32'd63; 
32'd1958: dataIn2 = 32'd59; 
32'd1959: dataIn2 = 32'd8; 
32'd1960: dataIn2 = 32'd90; 
32'd1961: dataIn2 = 32'd68; 
32'd1962: dataIn2 = 32'd98; 
32'd1963: dataIn2 = 32'd55; 
32'd1964: dataIn2 = 32'd52; 
32'd1965: dataIn2 = 32'd52; 
32'd1966: dataIn2 = 32'd100; 
32'd1967: dataIn2 = 32'd89; 
32'd1968: dataIn2 = 32'd56; 
32'd1969: dataIn2 = 32'd94; 
32'd1970: dataIn2 = 32'd73; 
32'd1971: dataIn2 = 32'd61; 
32'd1972: dataIn2 = 32'd51; 
32'd1973: dataIn2 = 32'd97; 
32'd1974: dataIn2 = 32'd48; 
32'd1975: dataIn2 = 32'd29; 
32'd1976: dataIn2 = 32'd91; 
32'd1977: dataIn2 = 32'd85; 
32'd1978: dataIn2 = 32'd58; 
32'd1979: dataIn2 = 32'd66; 
32'd1980: dataIn2 = 32'd4; 
32'd1981: dataIn2 = 32'd88; 
32'd1982: dataIn2 = 32'd55; 
32'd1983: dataIn2 = 32'd41; 
32'd1984: dataIn2 = 32'd11; 
32'd1985: dataIn2 = 32'd6; 
32'd1986: dataIn2 = 32'd81; 
32'd1987: dataIn2 = 32'd14; 
32'd1988: dataIn2 = 32'd36; 
32'd1989: dataIn2 = 32'd42; 
32'd1990: dataIn2 = 32'd17; 
32'd1991: dataIn2 = 32'd31; 
32'd1992: dataIn2 = 32'd27; 
32'd1993: dataIn2 = 32'd20; 
32'd1994: dataIn2 = 32'd5; 
32'd1995: dataIn2 = 32'd82; 
32'd1996: dataIn2 = 32'd4; 
32'd1997: dataIn2 = 32'd23; 
32'd1998: dataIn2 = 32'd27; 
32'd1999: dataIn2 = 32'd27; 
32'd2000: dataIn2 = 32'd39; 
32'd2001: dataIn2 = 32'd43; 
32'd2002: dataIn2 = 32'd62; 
32'd2003: dataIn2 = 32'd45; 
32'd2004: dataIn2 = 32'd15; 
32'd2005: dataIn2 = 32'd29; 
32'd2006: dataIn2 = 32'd98; 
32'd2007: dataIn2 = 32'd33; 
32'd2008: dataIn2 = 32'd98; 
32'd2009: dataIn2 = 32'd19; 
32'd2010: dataIn2 = 32'd99; 
32'd2011: dataIn2 = 32'd55; 
32'd2012: dataIn2 = 32'd88; 
32'd2013: dataIn2 = 32'd26; 
32'd2014: dataIn2 = 32'd64; 
32'd2015: dataIn2 = 32'd40; 
32'd2016: dataIn2 = 32'd36; 
32'd2017: dataIn2 = 32'd21; 
32'd2018: dataIn2 = 32'd38; 
32'd2019: dataIn2 = 32'd22; 
32'd2020: dataIn2 = 32'd81; 
32'd2021: dataIn2 = 32'd63; 
32'd2022: dataIn2 = 32'd17; 
32'd2023: dataIn2 = 32'd69; 
32'd2024: dataIn2 = 32'd46; 
32'd2025: dataIn2 = 32'd1; 
32'd2026: dataIn2 = 32'd27; 
32'd2027: dataIn2 = 32'd23; 
32'd2028: dataIn2 = 32'd74; 
32'd2029: dataIn2 = 32'd26; 
32'd2030: dataIn2 = 32'd84; 
32'd2031: dataIn2 = 32'd99; 
32'd2032: dataIn2 = 32'd100; 
32'd2033: dataIn2 = 32'd46; 
32'd2034: dataIn2 = 32'd30; 
32'd2035: dataIn2 = 32'd27; 
32'd2036: dataIn2 = 32'd85; 
32'd2037: dataIn2 = 32'd64; 
32'd2038: dataIn2 = 32'd15; 
32'd2039: dataIn2 = 32'd84; 
32'd2040: dataIn2 = 32'd92; 
32'd2041: dataIn2 = 32'd72; 
32'd2042: dataIn2 = 32'd69; 
32'd2043: dataIn2 = 32'd19; 
32'd2044: dataIn2 = 32'd79; 
32'd2045: dataIn2 = 32'd52; 
32'd2046: dataIn2 = 32'd100; 
32'd2047: dataIn2 = 32'd86; 
32'd2048: dataIn2 = 32'd96; 
32'd2049: dataIn2 = 32'd81; 
32'd2050: dataIn2 = 32'd58; 
32'd2051: dataIn2 = 32'd57; 
32'd2052: dataIn2 = 32'd84; 
32'd2053: dataIn2 = 32'd77; 
32'd2054: dataIn2 = 32'd66; 
32'd2055: dataIn2 = 32'd30; 
32'd2056: dataIn2 = 32'd36; 
32'd2057: dataIn2 = 32'd81; 
32'd2058: dataIn2 = 32'd38; 
32'd2059: dataIn2 = 32'd48; 
32'd2060: dataIn2 = 32'd95; 
32'd2061: dataIn2 = 32'd85; 
32'd2062: dataIn2 = 32'd43; 
32'd2063: dataIn2 = 32'd90; 
32'd2064: dataIn2 = 32'd16; 
32'd2065: dataIn2 = 32'd56; 
32'd2066: dataIn2 = 32'd49; 
32'd2067: dataIn2 = 32'd49; 
32'd2068: dataIn2 = 32'd28; 
32'd2069: dataIn2 = 32'd81; 
32'd2070: dataIn2 = 32'd0; 
32'd2071: dataIn2 = 32'd94; 
32'd2072: dataIn2 = 32'd83; 
32'd2073: dataIn2 = 32'd48; 
32'd2074: dataIn2 = 32'd88; 
32'd2075: dataIn2 = 32'd85; 
32'd2076: dataIn2 = 32'd87; 
32'd2077: dataIn2 = 32'd18; 
32'd2078: dataIn2 = 32'd86; 
32'd2079: dataIn2 = 32'd8; 
32'd2080: dataIn2 = 32'd77; 
32'd2081: dataIn2 = 32'd57; 
32'd2082: dataIn2 = 32'd4; 
32'd2083: dataIn2 = 32'd39; 
32'd2084: dataIn2 = 32'd76; 
32'd2085: dataIn2 = 32'd93; 
32'd2086: dataIn2 = 32'd44; 
32'd2087: dataIn2 = 32'd5; 
32'd2088: dataIn2 = 32'd84; 
32'd2089: dataIn2 = 32'd21; 
32'd2090: dataIn2 = 32'd75; 
32'd2091: dataIn2 = 32'd74; 
32'd2092: dataIn2 = 32'd68; 
32'd2093: dataIn2 = 32'd83; 
32'd2094: dataIn2 = 32'd9; 
32'd2095: dataIn2 = 32'd67; 
32'd2096: dataIn2 = 32'd98; 
32'd2097: dataIn2 = 32'd45; 
32'd2098: dataIn2 = 32'd93; 
32'd2099: dataIn2 = 32'd4; 
32'd2100: dataIn2 = 32'd55; 
32'd2101: dataIn2 = 32'd74; 
32'd2102: dataIn2 = 32'd24; 
32'd2103: dataIn2 = 32'd83; 
32'd2104: dataIn2 = 32'd70; 
32'd2105: dataIn2 = 32'd34; 
32'd2106: dataIn2 = 32'd18; 
32'd2107: dataIn2 = 32'd99; 
32'd2108: dataIn2 = 32'd53; 
32'd2109: dataIn2 = 32'd88; 
32'd2110: dataIn2 = 32'd64; 
32'd2111: dataIn2 = 32'd26; 
32'd2112: dataIn2 = 32'd40; 
32'd2113: dataIn2 = 32'd73; 
32'd2114: dataIn2 = 32'd38; 
32'd2115: dataIn2 = 32'd76; 
32'd2116: dataIn2 = 32'd77; 
32'd2117: dataIn2 = 32'd34; 
32'd2118: dataIn2 = 32'd49; 
32'd2119: dataIn2 = 32'd83; 
32'd2120: dataIn2 = 32'd9; 
32'd2121: dataIn2 = 32'd86; 
32'd2122: dataIn2 = 32'd47; 
32'd2123: dataIn2 = 32'd21; 
32'd2124: dataIn2 = 32'd80; 
32'd2125: dataIn2 = 32'd3; 
32'd2126: dataIn2 = 32'd42; 
32'd2127: dataIn2 = 32'd5; 
32'd2128: dataIn2 = 32'd32; 
32'd2129: dataIn2 = 32'd59; 
32'd2130: dataIn2 = 32'd46; 
32'd2131: dataIn2 = 32'd73; 
32'd2132: dataIn2 = 32'd48; 
32'd2133: dataIn2 = 32'd24; 
32'd2134: dataIn2 = 32'd60; 
32'd2135: dataIn2 = 32'd17; 
32'd2136: dataIn2 = 32'd17; 
32'd2137: dataIn2 = 32'd84; 
32'd2138: dataIn2 = 32'd66; 
32'd2139: dataIn2 = 32'd0; 
32'd2140: dataIn2 = 32'd32; 
32'd2141: dataIn2 = 32'd83; 
32'd2142: dataIn2 = 32'd37; 
32'd2143: dataIn2 = 32'd80; 
32'd2144: dataIn2 = 32'd8; 
32'd2145: dataIn2 = 32'd61; 
32'd2146: dataIn2 = 32'd30; 
32'd2147: dataIn2 = 32'd95; 
32'd2148: dataIn2 = 32'd98; 
32'd2149: dataIn2 = 32'd11; 
32'd2150: dataIn2 = 32'd42; 
32'd2151: dataIn2 = 32'd72; 
32'd2152: dataIn2 = 32'd87; 
32'd2153: dataIn2 = 32'd73; 
32'd2154: dataIn2 = 32'd57; 
32'd2155: dataIn2 = 32'd57; 
32'd2156: dataIn2 = 32'd18; 
32'd2157: dataIn2 = 32'd78; 
32'd2158: dataIn2 = 32'd29; 
32'd2159: dataIn2 = 32'd49; 
32'd2160: dataIn2 = 32'd66; 
32'd2161: dataIn2 = 32'd57; 
32'd2162: dataIn2 = 32'd28; 
32'd2163: dataIn2 = 32'd96; 
32'd2164: dataIn2 = 32'd58; 
32'd2165: dataIn2 = 32'd22; 
32'd2166: dataIn2 = 32'd89; 
32'd2167: dataIn2 = 32'd37; 
32'd2168: dataIn2 = 32'd43; 
32'd2169: dataIn2 = 32'd72; 
32'd2170: dataIn2 = 32'd43; 
32'd2171: dataIn2 = 32'd64; 
32'd2172: dataIn2 = 32'd25; 
32'd2173: dataIn2 = 32'd46; 
32'd2174: dataIn2 = 32'd17; 
32'd2175: dataIn2 = 32'd33; 
32'd2176: dataIn2 = 32'd50; 
32'd2177: dataIn2 = 32'd100; 
32'd2178: dataIn2 = 32'd32; 
32'd2179: dataIn2 = 32'd1; 
32'd2180: dataIn2 = 32'd70; 
32'd2181: dataIn2 = 32'd9; 
32'd2182: dataIn2 = 32'd86; 
32'd2183: dataIn2 = 32'd20; 
32'd2184: dataIn2 = 32'd94; 
32'd2185: dataIn2 = 32'd87; 
32'd2186: dataIn2 = 32'd47; 
32'd2187: dataIn2 = 32'd53; 
32'd2188: dataIn2 = 32'd94; 
32'd2189: dataIn2 = 32'd23; 
32'd2190: dataIn2 = 32'd91; 
32'd2191: dataIn2 = 32'd89; 
32'd2192: dataIn2 = 32'd77; 
32'd2193: dataIn2 = 32'd89; 
32'd2194: dataIn2 = 32'd24; 
32'd2195: dataIn2 = 32'd41; 
32'd2196: dataIn2 = 32'd11; 
32'd2197: dataIn2 = 32'd99; 
32'd2198: dataIn2 = 32'd83; 
32'd2199: dataIn2 = 32'd5; 
32'd2200: dataIn2 = 32'd54; 
32'd2201: dataIn2 = 32'd71; 
32'd2202: dataIn2 = 32'd95; 
32'd2203: dataIn2 = 32'd64; 
32'd2204: dataIn2 = 32'd86; 
32'd2205: dataIn2 = 32'd49; 
32'd2206: dataIn2 = 32'd96; 
32'd2207: dataIn2 = 32'd32; 
32'd2208: dataIn2 = 32'd92; 
32'd2209: dataIn2 = 32'd44; 
32'd2210: dataIn2 = 32'd37; 
32'd2211: dataIn2 = 32'd42; 
32'd2212: dataIn2 = 32'd12; 
32'd2213: dataIn2 = 32'd50; 
32'd2214: dataIn2 = 32'd83; 
32'd2215: dataIn2 = 32'd57; 
32'd2216: dataIn2 = 32'd33; 
32'd2217: dataIn2 = 32'd5; 
32'd2218: dataIn2 = 32'd42; 
32'd2219: dataIn2 = 32'd80; 
32'd2220: dataIn2 = 32'd38; 
32'd2221: dataIn2 = 32'd14; 
32'd2222: dataIn2 = 32'd63; 
32'd2223: dataIn2 = 32'd70; 
32'd2224: dataIn2 = 32'd67; 
32'd2225: dataIn2 = 32'd97; 
32'd2226: dataIn2 = 32'd69; 
32'd2227: dataIn2 = 32'd82; 
32'd2228: dataIn2 = 32'd73; 
32'd2229: dataIn2 = 32'd69; 
32'd2230: dataIn2 = 32'd12; 
32'd2231: dataIn2 = 32'd67; 
32'd2232: dataIn2 = 32'd99; 
32'd2233: dataIn2 = 32'd58; 
32'd2234: dataIn2 = 32'd71; 
32'd2235: dataIn2 = 32'd93; 
32'd2236: dataIn2 = 32'd13; 
32'd2237: dataIn2 = 32'd51; 
32'd2238: dataIn2 = 32'd55; 
32'd2239: dataIn2 = 32'd5; 
32'd2240: dataIn2 = 32'd86; 
32'd2241: dataIn2 = 32'd3; 
32'd2242: dataIn2 = 32'd64; 
32'd2243: dataIn2 = 32'd78; 
32'd2244: dataIn2 = 32'd36; 
32'd2245: dataIn2 = 32'd91; 
32'd2246: dataIn2 = 32'd94; 
32'd2247: dataIn2 = 32'd12; 
32'd2248: dataIn2 = 32'd31; 
32'd2249: dataIn2 = 32'd72; 
32'd2250: dataIn2 = 32'd61; 
32'd2251: dataIn2 = 32'd66; 
32'd2252: dataIn2 = 32'd99; 
32'd2253: dataIn2 = 32'd83; 
32'd2254: dataIn2 = 32'd90; 
32'd2255: dataIn2 = 32'd5; 
32'd2256: dataIn2 = 32'd46; 
32'd2257: dataIn2 = 32'd47; 
32'd2258: dataIn2 = 32'd68; 
32'd2259: dataIn2 = 32'd33; 
32'd2260: dataIn2 = 32'd34; 
32'd2261: dataIn2 = 32'd94; 
32'd2262: dataIn2 = 32'd57; 
32'd2263: dataIn2 = 32'd82; 
32'd2264: dataIn2 = 32'd3; 
32'd2265: dataIn2 = 32'd26; 
32'd2266: dataIn2 = 32'd85; 
32'd2267: dataIn2 = 32'd52; 
32'd2268: dataIn2 = 32'd88; 
32'd2269: dataIn2 = 32'd2; 
32'd2270: dataIn2 = 32'd55; 
32'd2271: dataIn2 = 32'd93; 
32'd2272: dataIn2 = 32'd65; 
32'd2273: dataIn2 = 32'd99; 
32'd2274: dataIn2 = 32'd30; 
32'd2275: dataIn2 = 32'd2; 
32'd2276: dataIn2 = 32'd95; 
32'd2277: dataIn2 = 32'd0; 
32'd2278: dataIn2 = 32'd36; 
32'd2279: dataIn2 = 32'd53; 
32'd2280: dataIn2 = 32'd89; 
32'd2281: dataIn2 = 32'd44; 
32'd2282: dataIn2 = 32'd69; 
32'd2283: dataIn2 = 32'd16; 
32'd2284: dataIn2 = 32'd9; 
32'd2285: dataIn2 = 32'd97; 
32'd2286: dataIn2 = 32'd21; 
32'd2287: dataIn2 = 32'd41; 
32'd2288: dataIn2 = 32'd44; 
32'd2289: dataIn2 = 32'd63; 
32'd2290: dataIn2 = 32'd73; 
32'd2291: dataIn2 = 32'd98; 
32'd2292: dataIn2 = 32'd23; 
32'd2293: dataIn2 = 32'd38; 
32'd2294: dataIn2 = 32'd73; 
32'd2295: dataIn2 = 32'd89; 
32'd2296: dataIn2 = 32'd87; 
32'd2297: dataIn2 = 32'd27; 
32'd2298: dataIn2 = 32'd86; 
32'd2299: dataIn2 = 32'd90; 
32'd2300: dataIn2 = 32'd6; 
32'd2301: dataIn2 = 32'd46; 
32'd2302: dataIn2 = 32'd11; 
32'd2303: dataIn2 = 32'd53; 
32'd2304: dataIn2 = 32'd33; 
32'd2305: dataIn2 = 32'd68; 
32'd2306: dataIn2 = 32'd58; 
32'd2307: dataIn2 = 32'd21; 
32'd2308: dataIn2 = 32'd90; 
32'd2309: dataIn2 = 32'd53; 
32'd2310: dataIn2 = 32'd16; 
32'd2311: dataIn2 = 32'd7; 
32'd2312: dataIn2 = 32'd88; 
32'd2313: dataIn2 = 32'd26; 
32'd2314: dataIn2 = 32'd20; 
32'd2315: dataIn2 = 32'd26; 
32'd2316: dataIn2 = 32'd89; 
32'd2317: dataIn2 = 32'd52; 
32'd2318: dataIn2 = 32'd5; 
32'd2319: dataIn2 = 32'd21; 
32'd2320: dataIn2 = 32'd91; 
32'd2321: dataIn2 = 32'd74; 
32'd2322: dataIn2 = 32'd12; 
32'd2323: dataIn2 = 32'd83; 
32'd2324: dataIn2 = 32'd50; 
32'd2325: dataIn2 = 32'd99; 
32'd2326: dataIn2 = 32'd49; 
32'd2327: dataIn2 = 32'd37; 
32'd2328: dataIn2 = 32'd45; 
32'd2329: dataIn2 = 32'd57; 
32'd2330: dataIn2 = 32'd90; 
32'd2331: dataIn2 = 32'd8; 
32'd2332: dataIn2 = 32'd70; 
32'd2333: dataIn2 = 32'd26; 
32'd2334: dataIn2 = 32'd82; 
32'd2335: dataIn2 = 32'd3; 
32'd2336: dataIn2 = 32'd12; 
32'd2337: dataIn2 = 32'd78; 
32'd2338: dataIn2 = 32'd61; 
32'd2339: dataIn2 = 32'd44; 
32'd2340: dataIn2 = 32'd36; 
32'd2341: dataIn2 = 32'd55; 
32'd2342: dataIn2 = 32'd35; 
32'd2343: dataIn2 = 32'd74; 
32'd2344: dataIn2 = 32'd19; 
32'd2345: dataIn2 = 32'd79; 
32'd2346: dataIn2 = 32'd44; 
32'd2347: dataIn2 = 32'd92; 
32'd2348: dataIn2 = 32'd33; 
32'd2349: dataIn2 = 32'd20; 
32'd2350: dataIn2 = 32'd50; 
32'd2351: dataIn2 = 32'd13; 
32'd2352: dataIn2 = 32'd28; 
32'd2353: dataIn2 = 32'd44; 
32'd2354: dataIn2 = 32'd23; 
32'd2355: dataIn2 = 32'd75; 
32'd2356: dataIn2 = 32'd4; 
32'd2357: dataIn2 = 32'd94; 
32'd2358: dataIn2 = 32'd35; 
32'd2359: dataIn2 = 32'd12; 
32'd2360: dataIn2 = 32'd26; 
32'd2361: dataIn2 = 32'd53; 
32'd2362: dataIn2 = 32'd93; 
32'd2363: dataIn2 = 32'd23; 
32'd2364: dataIn2 = 32'd80; 
32'd2365: dataIn2 = 32'd31; 
32'd2366: dataIn2 = 32'd98; 
32'd2367: dataIn2 = 32'd16; 
32'd2368: dataIn2 = 32'd98; 
32'd2369: dataIn2 = 32'd34; 
32'd2370: dataIn2 = 32'd92; 
32'd2371: dataIn2 = 32'd76; 
32'd2372: dataIn2 = 32'd55; 
32'd2373: dataIn2 = 32'd64; 
32'd2374: dataIn2 = 32'd26; 
32'd2375: dataIn2 = 32'd67; 
32'd2376: dataIn2 = 32'd74; 
32'd2377: dataIn2 = 32'd58; 
32'd2378: dataIn2 = 32'd21; 
32'd2379: dataIn2 = 32'd69; 
32'd2380: dataIn2 = 32'd37; 
32'd2381: dataIn2 = 32'd10; 
32'd2382: dataIn2 = 32'd83; 
32'd2383: dataIn2 = 32'd25; 
32'd2384: dataIn2 = 32'd72; 
32'd2385: dataIn2 = 32'd0; 
32'd2386: dataIn2 = 32'd74; 
32'd2387: dataIn2 = 32'd78; 
32'd2388: dataIn2 = 32'd66; 
32'd2389: dataIn2 = 32'd38; 
32'd2390: dataIn2 = 32'd85; 
32'd2391: dataIn2 = 32'd82; 
32'd2392: dataIn2 = 32'd23; 
32'd2393: dataIn2 = 32'd17; 
32'd2394: dataIn2 = 32'd12; 
32'd2395: dataIn2 = 32'd92; 
32'd2396: dataIn2 = 32'd10; 
32'd2397: dataIn2 = 32'd15; 
32'd2398: dataIn2 = 32'd49; 
32'd2399: dataIn2 = 32'd25; 
32'd2400: dataIn2 = 32'd12; 
32'd2401: dataIn2 = 32'd68; 
32'd2402: dataIn2 = 32'd18; 
32'd2403: dataIn2 = 32'd88; 
32'd2404: dataIn2 = 32'd2; 
32'd2405: dataIn2 = 32'd80; 
32'd2406: dataIn2 = 32'd100; 
32'd2407: dataIn2 = 32'd27; 
32'd2408: dataIn2 = 32'd44; 
32'd2409: dataIn2 = 32'd16; 
32'd2410: dataIn2 = 32'd50; 
32'd2411: dataIn2 = 32'd49; 
32'd2412: dataIn2 = 32'd39; 
32'd2413: dataIn2 = 32'd0; 
32'd2414: dataIn2 = 32'd53; 
32'd2415: dataIn2 = 32'd100; 
32'd2416: dataIn2 = 32'd52; 
32'd2417: dataIn2 = 32'd5; 
32'd2418: dataIn2 = 32'd76; 
32'd2419: dataIn2 = 32'd71; 
32'd2420: dataIn2 = 32'd55; 
32'd2421: dataIn2 = 32'd43; 
32'd2422: dataIn2 = 32'd31; 
32'd2423: dataIn2 = 32'd35; 
32'd2424: dataIn2 = 32'd84; 
32'd2425: dataIn2 = 32'd28; 
32'd2426: dataIn2 = 32'd46; 
32'd2427: dataIn2 = 32'd47; 
32'd2428: dataIn2 = 32'd46; 
32'd2429: dataIn2 = 32'd83; 
32'd2430: dataIn2 = 32'd25; 
32'd2431: dataIn2 = 32'd76; 
32'd2432: dataIn2 = 32'd49; 
32'd2433: dataIn2 = 32'd61; 
32'd2434: dataIn2 = 32'd19; 
32'd2435: dataIn2 = 32'd94; 
32'd2436: dataIn2 = 32'd74; 
32'd2437: dataIn2 = 32'd56; 
32'd2438: dataIn2 = 32'd95; 
32'd2439: dataIn2 = 32'd80; 
32'd2440: dataIn2 = 32'd62; 
32'd2441: dataIn2 = 32'd84; 
32'd2442: dataIn2 = 32'd38; 
32'd2443: dataIn2 = 32'd94; 
32'd2444: dataIn2 = 32'd14; 
32'd2445: dataIn2 = 32'd9; 
32'd2446: dataIn2 = 32'd41; 
32'd2447: dataIn2 = 32'd13; 
32'd2448: dataIn2 = 32'd59; 
32'd2449: dataIn2 = 32'd93; 
32'd2450: dataIn2 = 32'd78; 
32'd2451: dataIn2 = 32'd93; 
32'd2452: dataIn2 = 32'd55; 
32'd2453: dataIn2 = 32'd15; 
32'd2454: dataIn2 = 32'd88; 
32'd2455: dataIn2 = 32'd38; 
32'd2456: dataIn2 = 32'd68; 
32'd2457: dataIn2 = 32'd65; 
32'd2458: dataIn2 = 32'd10; 
32'd2459: dataIn2 = 32'd68; 
32'd2460: dataIn2 = 32'd56; 
32'd2461: dataIn2 = 32'd55; 
32'd2462: dataIn2 = 32'd71; 
32'd2463: dataIn2 = 32'd5; 
32'd2464: dataIn2 = 32'd90; 
32'd2465: dataIn2 = 32'd83; 
32'd2466: dataIn2 = 32'd3; 
32'd2467: dataIn2 = 32'd48; 
32'd2468: dataIn2 = 32'd39; 
32'd2469: dataIn2 = 32'd17; 
32'd2470: dataIn2 = 32'd92; 
32'd2471: dataIn2 = 32'd37; 
32'd2472: dataIn2 = 32'd95; 
32'd2473: dataIn2 = 32'd43; 
32'd2474: dataIn2 = 32'd93; 
32'd2475: dataIn2 = 32'd47; 
32'd2476: dataIn2 = 32'd53; 
32'd2477: dataIn2 = 32'd22; 
32'd2478: dataIn2 = 32'd5; 
32'd2479: dataIn2 = 32'd28; 
32'd2480: dataIn2 = 32'd24; 
32'd2481: dataIn2 = 32'd69; 
32'd2482: dataIn2 = 32'd61; 
32'd2483: dataIn2 = 32'd5; 
32'd2484: dataIn2 = 32'd46; 
32'd2485: dataIn2 = 32'd88; 
32'd2486: dataIn2 = 32'd51; 
32'd2487: dataIn2 = 32'd9; 
32'd2488: dataIn2 = 32'd72; 
32'd2489: dataIn2 = 32'd75; 
32'd2490: dataIn2 = 32'd58; 
32'd2491: dataIn2 = 32'd35; 
32'd2492: dataIn2 = 32'd87; 
32'd2493: dataIn2 = 32'd38; 
32'd2494: dataIn2 = 32'd55; 
32'd2495: dataIn2 = 32'd25; 
32'd2496: dataIn2 = 32'd19; 
32'd2497: dataIn2 = 32'd20; 
32'd2498: dataIn2 = 32'd73; 
32'd2499: dataIn2 = 32'd26; 
32'd2500: dataIn2 = 32'd3; 
32'd2501: dataIn2 = 32'd70; 
32'd2502: dataIn2 = 32'd90; 
32'd2503: dataIn2 = 32'd93; 
32'd2504: dataIn2 = 32'd27; 
32'd2505: dataIn2 = 32'd64; 
32'd2506: dataIn2 = 32'd70; 
32'd2507: dataIn2 = 32'd66; 
32'd2508: dataIn2 = 32'd35; 
32'd2509: dataIn2 = 32'd73; 
32'd2510: dataIn2 = 32'd55; 
32'd2511: dataIn2 = 32'd23; 
32'd2512: dataIn2 = 32'd65; 
32'd2513: dataIn2 = 32'd19; 
32'd2514: dataIn2 = 32'd2; 
32'd2515: dataIn2 = 32'd6; 
32'd2516: dataIn2 = 32'd77; 
32'd2517: dataIn2 = 32'd67; 
32'd2518: dataIn2 = 32'd46; 
32'd2519: dataIn2 = 32'd69; 
32'd2520: dataIn2 = 32'd73; 
32'd2521: dataIn2 = 32'd85; 
32'd2522: dataIn2 = 32'd70; 
32'd2523: dataIn2 = 32'd39; 
32'd2524: dataIn2 = 32'd88; 
32'd2525: dataIn2 = 32'd60; 
32'd2526: dataIn2 = 32'd6; 
32'd2527: dataIn2 = 32'd62; 
32'd2528: dataIn2 = 32'd22; 
32'd2529: dataIn2 = 32'd17; 
32'd2530: dataIn2 = 32'd14; 
32'd2531: dataIn2 = 32'd34; 
32'd2532: dataIn2 = 32'd48; 
32'd2533: dataIn2 = 32'd17; 
32'd2534: dataIn2 = 32'd32; 
32'd2535: dataIn2 = 32'd0; 
32'd2536: dataIn2 = 32'd84; 
32'd2537: dataIn2 = 32'd1; 
32'd2538: dataIn2 = 32'd23; 
32'd2539: dataIn2 = 32'd26; 
32'd2540: dataIn2 = 32'd38; 
32'd2541: dataIn2 = 32'd68; 
32'd2542: dataIn2 = 32'd19; 
32'd2543: dataIn2 = 32'd21; 
32'd2544: dataIn2 = 32'd95; 
32'd2545: dataIn2 = 32'd98; 
32'd2546: dataIn2 = 32'd55; 
32'd2547: dataIn2 = 32'd19; 
32'd2548: dataIn2 = 32'd14; 
32'd2549: dataIn2 = 32'd13; 
32'd2550: dataIn2 = 32'd71; 
32'd2551: dataIn2 = 32'd89; 
32'd2552: dataIn2 = 32'd84; 
32'd2553: dataIn2 = 32'd43; 
32'd2554: dataIn2 = 32'd13; 
32'd2555: dataIn2 = 32'd51; 
32'd2556: dataIn2 = 32'd18; 
32'd2557: dataIn2 = 32'd88; 
32'd2558: dataIn2 = 32'd45; 
32'd2559: dataIn2 = 32'd0; 
32'd2560: dataIn2 = 32'd5; 
32'd2561: dataIn2 = 32'd53; 
32'd2562: dataIn2 = 32'd61; 
32'd2563: dataIn2 = 32'd13; 
32'd2564: dataIn2 = 32'd97; 
32'd2565: dataIn2 = 32'd59; 
32'd2566: dataIn2 = 32'd45; 
32'd2567: dataIn2 = 32'd4; 
32'd2568: dataIn2 = 32'd92; 
32'd2569: dataIn2 = 32'd44; 
32'd2570: dataIn2 = 32'd35; 
32'd2571: dataIn2 = 32'd0; 
32'd2572: dataIn2 = 32'd35; 
32'd2573: dataIn2 = 32'd62; 
32'd2574: dataIn2 = 32'd20; 
32'd2575: dataIn2 = 32'd15; 
32'd2576: dataIn2 = 32'd46; 
32'd2577: dataIn2 = 32'd45; 
32'd2578: dataIn2 = 32'd5; 
32'd2579: dataIn2 = 32'd36; 
32'd2580: dataIn2 = 32'd67; 
32'd2581: dataIn2 = 32'd90; 
32'd2582: dataIn2 = 32'd17; 
32'd2583: dataIn2 = 32'd61; 
32'd2584: dataIn2 = 32'd97; 
32'd2585: dataIn2 = 32'd5; 
32'd2586: dataIn2 = 32'd78; 
32'd2587: dataIn2 = 32'd77; 
32'd2588: dataIn2 = 32'd65; 
32'd2589: dataIn2 = 32'd86; 
32'd2590: dataIn2 = 32'd80; 
32'd2591: dataIn2 = 32'd39; 
32'd2592: dataIn2 = 32'd93; 
32'd2593: dataIn2 = 32'd100; 
32'd2594: dataIn2 = 32'd96; 
32'd2595: dataIn2 = 32'd11; 
32'd2596: dataIn2 = 32'd74; 
32'd2597: dataIn2 = 32'd39; 
32'd2598: dataIn2 = 32'd28; 
32'd2599: dataIn2 = 32'd71; 
32'd2600: dataIn2 = 32'd46; 
32'd2601: dataIn2 = 32'd87; 
32'd2602: dataIn2 = 32'd4; 
32'd2603: dataIn2 = 32'd42; 
32'd2604: dataIn2 = 32'd48; 
32'd2605: dataIn2 = 32'd14; 
32'd2606: dataIn2 = 32'd11; 
32'd2607: dataIn2 = 32'd2; 
32'd2608: dataIn2 = 32'd53; 
32'd2609: dataIn2 = 32'd12; 
32'd2610: dataIn2 = 32'd27; 
32'd2611: dataIn2 = 32'd4; 
32'd2612: dataIn2 = 32'd97; 
32'd2613: dataIn2 = 32'd83; 
32'd2614: dataIn2 = 32'd18; 
32'd2615: dataIn2 = 32'd32; 
32'd2616: dataIn2 = 32'd50; 
32'd2617: dataIn2 = 32'd63; 
32'd2618: dataIn2 = 32'd42; 
32'd2619: dataIn2 = 32'd18; 
32'd2620: dataIn2 = 32'd61; 
32'd2621: dataIn2 = 32'd36; 
32'd2622: dataIn2 = 32'd74; 
32'd2623: dataIn2 = 32'd80; 
32'd2624: dataIn2 = 32'd14; 
32'd2625: dataIn2 = 32'd32; 
32'd2626: dataIn2 = 32'd44; 
32'd2627: dataIn2 = 32'd8; 
32'd2628: dataIn2 = 32'd58; 
32'd2629: dataIn2 = 32'd92; 
32'd2630: dataIn2 = 32'd94; 
32'd2631: dataIn2 = 32'd80; 
32'd2632: dataIn2 = 32'd54; 
32'd2633: dataIn2 = 32'd97; 
32'd2634: dataIn2 = 32'd89; 
32'd2635: dataIn2 = 32'd27; 
32'd2636: dataIn2 = 32'd73; 
32'd2637: dataIn2 = 32'd41; 
32'd2638: dataIn2 = 32'd90; 
32'd2639: dataIn2 = 32'd12; 
32'd2640: dataIn2 = 32'd28; 
32'd2641: dataIn2 = 32'd64; 
32'd2642: dataIn2 = 32'd68; 
32'd2643: dataIn2 = 32'd48; 
32'd2644: dataIn2 = 32'd33; 
32'd2645: dataIn2 = 32'd9; 
32'd2646: dataIn2 = 32'd62; 
32'd2647: dataIn2 = 32'd24; 
32'd2648: dataIn2 = 32'd15; 
32'd2649: dataIn2 = 32'd95; 
32'd2650: dataIn2 = 32'd29; 
32'd2651: dataIn2 = 32'd57; 
32'd2652: dataIn2 = 32'd3; 
32'd2653: dataIn2 = 32'd18; 
32'd2654: dataIn2 = 32'd94; 
32'd2655: dataIn2 = 32'd26; 
32'd2656: dataIn2 = 32'd58; 
32'd2657: dataIn2 = 32'd35; 
32'd2658: dataIn2 = 32'd92; 
32'd2659: dataIn2 = 32'd38; 
32'd2660: dataIn2 = 32'd50; 
32'd2661: dataIn2 = 32'd97; 
32'd2662: dataIn2 = 32'd54; 
32'd2663: dataIn2 = 32'd95; 
32'd2664: dataIn2 = 32'd36; 
32'd2665: dataIn2 = 32'd54; 
32'd2666: dataIn2 = 32'd62; 
32'd2667: dataIn2 = 32'd86; 
32'd2668: dataIn2 = 32'd87; 
32'd2669: dataIn2 = 32'd39; 
32'd2670: dataIn2 = 32'd21; 
32'd2671: dataIn2 = 32'd79; 
32'd2672: dataIn2 = 32'd34; 
32'd2673: dataIn2 = 32'd65; 
32'd2674: dataIn2 = 32'd10; 
32'd2675: dataIn2 = 32'd13; 
32'd2676: dataIn2 = 32'd64; 
32'd2677: dataIn2 = 32'd99; 
32'd2678: dataIn2 = 32'd0; 
32'd2679: dataIn2 = 32'd66; 
32'd2680: dataIn2 = 32'd43; 
32'd2681: dataIn2 = 32'd86; 
32'd2682: dataIn2 = 32'd13; 
32'd2683: dataIn2 = 32'd78; 
32'd2684: dataIn2 = 32'd96; 
32'd2685: dataIn2 = 32'd100; 
32'd2686: dataIn2 = 32'd14; 
32'd2687: dataIn2 = 32'd10; 
32'd2688: dataIn2 = 32'd20; 
32'd2689: dataIn2 = 32'd21; 
32'd2690: dataIn2 = 32'd48; 
32'd2691: dataIn2 = 32'd67; 
32'd2692: dataIn2 = 32'd84; 
32'd2693: dataIn2 = 32'd48; 
32'd2694: dataIn2 = 32'd30; 
32'd2695: dataIn2 = 32'd66; 
32'd2696: dataIn2 = 32'd25; 
32'd2697: dataIn2 = 32'd41; 
32'd2698: dataIn2 = 32'd55; 
32'd2699: dataIn2 = 32'd63; 
32'd2700: dataIn2 = 32'd35; 
32'd2701: dataIn2 = 32'd29; 
32'd2702: dataIn2 = 32'd4; 
32'd2703: dataIn2 = 32'd74; 
32'd2704: dataIn2 = 32'd18; 
32'd2705: dataIn2 = 32'd61; 
32'd2706: dataIn2 = 32'd5; 
32'd2707: dataIn2 = 32'd77; 
32'd2708: dataIn2 = 32'd83; 
32'd2709: dataIn2 = 32'd60; 
32'd2710: dataIn2 = 32'd67; 
32'd2711: dataIn2 = 32'd34; 
32'd2712: dataIn2 = 32'd58; 
32'd2713: dataIn2 = 32'd42; 
32'd2714: dataIn2 = 32'd76; 
32'd2715: dataIn2 = 32'd13; 
32'd2716: dataIn2 = 32'd89; 
32'd2717: dataIn2 = 32'd19; 
32'd2718: dataIn2 = 32'd0; 
32'd2719: dataIn2 = 32'd40; 
32'd2720: dataIn2 = 32'd14; 
32'd2721: dataIn2 = 32'd54; 
32'd2722: dataIn2 = 32'd87; 
32'd2723: dataIn2 = 32'd26; 
32'd2724: dataIn2 = 32'd50; 
32'd2725: dataIn2 = 32'd97; 
32'd2726: dataIn2 = 32'd69; 
32'd2727: dataIn2 = 32'd57; 
32'd2728: dataIn2 = 32'd2; 
32'd2729: dataIn2 = 32'd53; 
32'd2730: dataIn2 = 32'd66; 
32'd2731: dataIn2 = 32'd57; 
32'd2732: dataIn2 = 32'd1; 
32'd2733: dataIn2 = 32'd23; 
32'd2734: dataIn2 = 32'd21; 
32'd2735: dataIn2 = 32'd45; 
32'd2736: dataIn2 = 32'd62; 
32'd2737: dataIn2 = 32'd6; 
32'd2738: dataIn2 = 32'd2; 
32'd2739: dataIn2 = 32'd98; 
32'd2740: dataIn2 = 32'd88; 
32'd2741: dataIn2 = 32'd60; 
32'd2742: dataIn2 = 32'd71; 
32'd2743: dataIn2 = 32'd35; 
32'd2744: dataIn2 = 32'd43; 
32'd2745: dataIn2 = 32'd98; 
32'd2746: dataIn2 = 32'd82; 
32'd2747: dataIn2 = 32'd6; 
32'd2748: dataIn2 = 32'd35; 
32'd2749: dataIn2 = 32'd11; 
32'd2750: dataIn2 = 32'd32; 
32'd2751: dataIn2 = 32'd37; 
32'd2752: dataIn2 = 32'd23; 
32'd2753: dataIn2 = 32'd44; 
32'd2754: dataIn2 = 32'd23; 
32'd2755: dataIn2 = 32'd13; 
32'd2756: dataIn2 = 32'd71; 
32'd2757: dataIn2 = 32'd53; 
32'd2758: dataIn2 = 32'd23; 
32'd2759: dataIn2 = 32'd29; 
32'd2760: dataIn2 = 32'd45; 
32'd2761: dataIn2 = 32'd97; 
32'd2762: dataIn2 = 32'd62; 
32'd2763: dataIn2 = 32'd47; 
32'd2764: dataIn2 = 32'd49; 
32'd2765: dataIn2 = 32'd68; 
32'd2766: dataIn2 = 32'd29; 
32'd2767: dataIn2 = 32'd66; 
32'd2768: dataIn2 = 32'd2; 
32'd2769: dataIn2 = 32'd2; 
32'd2770: dataIn2 = 32'd83; 
32'd2771: dataIn2 = 32'd32; 
32'd2772: dataIn2 = 32'd80; 
32'd2773: dataIn2 = 32'd65; 
32'd2774: dataIn2 = 32'd67; 
32'd2775: dataIn2 = 32'd45; 
32'd2776: dataIn2 = 32'd36; 
32'd2777: dataIn2 = 32'd48; 
32'd2778: dataIn2 = 32'd16; 
32'd2779: dataIn2 = 32'd93; 
32'd2780: dataIn2 = 32'd84; 
32'd2781: dataIn2 = 32'd27; 
32'd2782: dataIn2 = 32'd10; 
32'd2783: dataIn2 = 32'd80; 
32'd2784: dataIn2 = 32'd30; 
32'd2785: dataIn2 = 32'd49; 
32'd2786: dataIn2 = 32'd71; 
32'd2787: dataIn2 = 32'd68; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_64_40.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
