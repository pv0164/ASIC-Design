//64x64 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 1229 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd330 ; 
  wdata_col_base = 32'd15590 ; 
  row_base = 32'd168190 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #138000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd168190: dataIn1 = 32'd0
; 
32'd168191: dataIn1 = 32'd20
; 
32'd168192: dataIn1 = 32'd40
; 
32'd168193: dataIn1 = 32'd54
; 
32'd168194: dataIn1 = 32'd74
; 
32'd168195: dataIn1 = 32'd100
; 
32'd168196: dataIn1 = 32'd117
; 
32'd168197: dataIn1 = 32'd136
; 
32'd168198: dataIn1 = 32'd156
; 
32'd168199: dataIn1 = 32'd173
; 
32'd168200: dataIn1 = 32'd191
; 
32'd168201: dataIn1 = 32'd208
; 
32'd168202: dataIn1 = 32'd217
; 
32'd168203: dataIn1 = 32'd238
; 
32'd168204: dataIn1 = 32'd256
; 
32'd168205: dataIn1 = 32'd276
; 
32'd168206: dataIn1 = 32'd297
; 
32'd168207: dataIn1 = 32'd313
; 
32'd168208: dataIn1 = 32'd334
; 
32'd168209: dataIn1 = 32'd354
; 
32'd168210: dataIn1 = 32'd378
; 
32'd168211: dataIn1 = 32'd399
; 
32'd168212: dataIn1 = 32'd421
; 
32'd168213: dataIn1 = 32'd436
; 
32'd168214: dataIn1 = 32'd454
; 
32'd168215: dataIn1 = 32'd482
; 
32'd168216: dataIn1 = 32'd498
; 
32'd168217: dataIn1 = 32'd518
; 
32'd168218: dataIn1 = 32'd536
; 
32'd168219: dataIn1 = 32'd551
; 
32'd168220: dataIn1 = 32'd569
; 
32'd168221: dataIn1 = 32'd588
; 
32'd168222: dataIn1 = 32'd603
; 
32'd168223: dataIn1 = 32'd623
; 
32'd168224: dataIn1 = 32'd637
; 
32'd168225: dataIn1 = 32'd655
; 
32'd168226: dataIn1 = 32'd672
; 
32'd168227: dataIn1 = 32'd693
; 
32'd168228: dataIn1 = 32'd707
; 
32'd168229: dataIn1 = 32'd724
; 
32'd168230: dataIn1 = 32'd740
; 
32'd168231: dataIn1 = 32'd761
; 
32'd168232: dataIn1 = 32'd776
; 
32'd168233: dataIn1 = 32'd799
; 
32'd168234: dataIn1 = 32'd817
; 
32'd168235: dataIn1 = 32'd840
; 
32'd168236: dataIn1 = 32'd855
; 
32'd168237: dataIn1 = 32'd880
; 
32'd168238: dataIn1 = 32'd899
; 
32'd168239: dataIn1 = 32'd916
; 
32'd168240: dataIn1 = 32'd934
; 
32'd168241: dataIn1 = 32'd946
; 
32'd168242: dataIn1 = 32'd962
; 
32'd168243: dataIn1 = 32'd985
; 
32'd168244: dataIn1 = 32'd1002
; 
32'd168245: dataIn1 = 32'd1029
; 
32'd168246: dataIn1 = 32'd1048
; 
32'd168247: dataIn1 = 32'd1068
; 
32'd168248: dataIn1 = 32'd1088
; 
32'd168249: dataIn1 = 32'd1110
; 
32'd168250: dataIn1 = 32'd1131
; 
32'd168251: dataIn1 = 32'd1147
; 
32'd168252: dataIn1 = 32'd1169
; 
32'd168253: dataIn1 = 32'd1189
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd15590: dataIn1 = 32'd0
; 
32'd15591: dataIn1 = 32'd20
; 
32'd15592: dataIn1 = 32'd40
; 
32'd15593: dataIn1 = 32'd54
; 
32'd15594: dataIn1 = 32'd74
; 
32'd15595: dataIn1 = 32'd100
; 
32'd15596: dataIn1 = 32'd117
; 
32'd15597: dataIn1 = 32'd136
; 
32'd15598: dataIn1 = 32'd156
; 
32'd15599: dataIn1 = 32'd173
; 
32'd15600: dataIn1 = 32'd191
; 
32'd15601: dataIn1 = 32'd208
; 
32'd15602: dataIn1 = 32'd217
; 
32'd15603: dataIn1 = 32'd238
; 
32'd15604: dataIn1 = 32'd256
; 
32'd15605: dataIn1 = 32'd276
; 
32'd15606: dataIn1 = 32'd297
; 
32'd15607: dataIn1 = 32'd313
; 
32'd15608: dataIn1 = 32'd334
; 
32'd15609: dataIn1 = 32'd354
; 
32'd15610: dataIn1 = 32'd378
; 
32'd15611: dataIn1 = 32'd399
; 
32'd15612: dataIn1 = 32'd421
; 
32'd15613: dataIn1 = 32'd436
; 
32'd15614: dataIn1 = 32'd454
; 
32'd15615: dataIn1 = 32'd482
; 
32'd15616: dataIn1 = 32'd498
; 
32'd15617: dataIn1 = 32'd518
; 
32'd15618: dataIn1 = 32'd536
; 
32'd15619: dataIn1 = 32'd551
; 
32'd15620: dataIn1 = 32'd569
; 
32'd15621: dataIn1 = 32'd588
; 
32'd15622: dataIn1 = 32'd603
; 
32'd15623: dataIn1 = 32'd623
; 
32'd15624: dataIn1 = 32'd637
; 
32'd15625: dataIn1 = 32'd655
; 
32'd15626: dataIn1 = 32'd672
; 
32'd15627: dataIn1 = 32'd693
; 
32'd15628: dataIn1 = 32'd707
; 
32'd15629: dataIn1 = 32'd724
; 
32'd15630: dataIn1 = 32'd740
; 
32'd15631: dataIn1 = 32'd761
; 
32'd15632: dataIn1 = 32'd776
; 
32'd15633: dataIn1 = 32'd799
; 
32'd15634: dataIn1 = 32'd817
; 
32'd15635: dataIn1 = 32'd840
; 
32'd15636: dataIn1 = 32'd855
; 
32'd15637: dataIn1 = 32'd880
; 
32'd15638: dataIn1 = 32'd899
; 
32'd15639: dataIn1 = 32'd916
; 
32'd15640: dataIn1 = 32'd934
; 
32'd15641: dataIn1 = 32'd946
; 
32'd15642: dataIn1 = 32'd962
; 
32'd15643: dataIn1 = 32'd985
; 
32'd15644: dataIn1 = 32'd1002
; 
32'd15645: dataIn1 = 32'd1029
; 
32'd15646: dataIn1 = 32'd1048
; 
32'd15647: dataIn1 = 32'd1068
; 
32'd15648: dataIn1 = 32'd1088
; 
32'd15649: dataIn1 = 32'd1110
; 
32'd15650: dataIn1 = 32'd1131
; 
32'd15651: dataIn1 = 32'd1147
; 
32'd15652: dataIn1 = 32'd1169
; 
32'd15653: dataIn1 = 32'd1189
; 
32'd15654: dataIn1 = 32'd1203
; 
32'd15655: dataIn1 = 32'd6
; 
32'd15656: dataIn1 = 32'd13
; 
32'd15657: dataIn1 = 32'd14
; 
32'd15658: dataIn1 = 32'd19
; 
32'd15659: dataIn1 = 32'd20
; 
32'd15660: dataIn1 = 32'd24
; 
32'd15661: dataIn1 = 32'd25
; 
32'd15662: dataIn1 = 32'd29
; 
32'd15663: dataIn1 = 32'd35
; 
32'd15664: dataIn1 = 32'd37
; 
32'd15665: dataIn1 = 32'd40
; 
32'd15666: dataIn1 = 32'd42
; 
32'd15667: dataIn1 = 32'd43
; 
32'd15668: dataIn1 = 32'd45
; 
32'd15669: dataIn1 = 32'd46
; 
32'd15670: dataIn1 = 32'd50
; 
32'd15671: dataIn1 = 32'd52
; 
32'd15672: dataIn1 = 32'd54
; 
32'd15673: dataIn1 = 32'd55
; 
32'd15674: dataIn1 = 32'd57
; 
32'd15675: dataIn1 = 32'd4
; 
32'd15676: dataIn1 = 32'd6
; 
32'd15677: dataIn1 = 32'd8
; 
32'd15678: dataIn1 = 32'd9
; 
32'd15679: dataIn1 = 32'd10
; 
32'd15680: dataIn1 = 32'd12
; 
32'd15681: dataIn1 = 32'd15
; 
32'd15682: dataIn1 = 32'd20
; 
32'd15683: dataIn1 = 32'd21
; 
32'd15684: dataIn1 = 32'd28
; 
32'd15685: dataIn1 = 32'd31
; 
32'd15686: dataIn1 = 32'd36
; 
32'd15687: dataIn1 = 32'd40
; 
32'd15688: dataIn1 = 32'd46
; 
32'd15689: dataIn1 = 32'd47
; 
32'd15690: dataIn1 = 32'd49
; 
32'd15691: dataIn1 = 32'd50
; 
32'd15692: dataIn1 = 32'd51
; 
32'd15693: dataIn1 = 32'd52
; 
32'd15694: dataIn1 = 32'd58
; 
32'd15695: dataIn1 = 32'd0
; 
32'd15696: dataIn1 = 32'd2
; 
32'd15697: dataIn1 = 32'd8
; 
32'd15698: dataIn1 = 32'd14
; 
32'd15699: dataIn1 = 32'd27
; 
32'd15700: dataIn1 = 32'd29
; 
32'd15701: dataIn1 = 32'd34
; 
32'd15702: dataIn1 = 32'd43
; 
32'd15703: dataIn1 = 32'd44
; 
32'd15704: dataIn1 = 32'd46
; 
32'd15705: dataIn1 = 32'd48
; 
32'd15706: dataIn1 = 32'd57
; 
32'd15707: dataIn1 = 32'd59
; 
32'd15708: dataIn1 = 32'd61
; 
32'd15709: dataIn1 = 32'd3
; 
32'd15710: dataIn1 = 32'd5
; 
32'd15711: dataIn1 = 32'd6
; 
32'd15712: dataIn1 = 32'd14
; 
32'd15713: dataIn1 = 32'd18
; 
32'd15714: dataIn1 = 32'd20
; 
32'd15715: dataIn1 = 32'd26
; 
32'd15716: dataIn1 = 32'd27
; 
32'd15717: dataIn1 = 32'd29
; 
32'd15718: dataIn1 = 32'd31
; 
32'd15719: dataIn1 = 32'd37
; 
32'd15720: dataIn1 = 32'd45
; 
32'd15721: dataIn1 = 32'd48
; 
32'd15722: dataIn1 = 32'd49
; 
32'd15723: dataIn1 = 32'd50
; 
32'd15724: dataIn1 = 32'd51
; 
32'd15725: dataIn1 = 32'd53
; 
32'd15726: dataIn1 = 32'd54
; 
32'd15727: dataIn1 = 32'd58
; 
32'd15728: dataIn1 = 32'd60
; 
32'd15729: dataIn1 = 32'd0
; 
32'd15730: dataIn1 = 32'd2
; 
32'd15731: dataIn1 = 32'd5
; 
32'd15732: dataIn1 = 32'd8
; 
32'd15733: dataIn1 = 32'd12
; 
32'd15734: dataIn1 = 32'd13
; 
32'd15735: dataIn1 = 32'd14
; 
32'd15736: dataIn1 = 32'd15
; 
32'd15737: dataIn1 = 32'd21
; 
32'd15738: dataIn1 = 32'd27
; 
32'd15739: dataIn1 = 32'd29
; 
32'd15740: dataIn1 = 32'd30
; 
32'd15741: dataIn1 = 32'd31
; 
32'd15742: dataIn1 = 32'd32
; 
32'd15743: dataIn1 = 32'd36
; 
32'd15744: dataIn1 = 32'd37
; 
32'd15745: dataIn1 = 32'd38
; 
32'd15746: dataIn1 = 32'd39
; 
32'd15747: dataIn1 = 32'd42
; 
32'd15748: dataIn1 = 32'd46
; 
32'd15749: dataIn1 = 32'd47
; 
32'd15750: dataIn1 = 32'd50
; 
32'd15751: dataIn1 = 32'd52
; 
32'd15752: dataIn1 = 32'd59
; 
32'd15753: dataIn1 = 32'd60
; 
32'd15754: dataIn1 = 32'd63
; 
32'd15755: dataIn1 = 32'd2
; 
32'd15756: dataIn1 = 32'd18
; 
32'd15757: dataIn1 = 32'd19
; 
32'd15758: dataIn1 = 32'd26
; 
32'd15759: dataIn1 = 32'd33
; 
32'd15760: dataIn1 = 32'd36
; 
32'd15761: dataIn1 = 32'd38
; 
32'd15762: dataIn1 = 32'd41
; 
32'd15763: dataIn1 = 32'd44
; 
32'd15764: dataIn1 = 32'd46
; 
32'd15765: dataIn1 = 32'd48
; 
32'd15766: dataIn1 = 32'd50
; 
32'd15767: dataIn1 = 32'd51
; 
32'd15768: dataIn1 = 32'd54
; 
32'd15769: dataIn1 = 32'd56
; 
32'd15770: dataIn1 = 32'd57
; 
32'd15771: dataIn1 = 32'd63
; 
32'd15772: dataIn1 = 32'd2
; 
32'd15773: dataIn1 = 32'd3
; 
32'd15774: dataIn1 = 32'd9
; 
32'd15775: dataIn1 = 32'd10
; 
32'd15776: dataIn1 = 32'd13
; 
32'd15777: dataIn1 = 32'd21
; 
32'd15778: dataIn1 = 32'd22
; 
32'd15779: dataIn1 = 32'd23
; 
32'd15780: dataIn1 = 32'd27
; 
32'd15781: dataIn1 = 32'd28
; 
32'd15782: dataIn1 = 32'd29
; 
32'd15783: dataIn1 = 32'd30
; 
32'd15784: dataIn1 = 32'd33
; 
32'd15785: dataIn1 = 32'd43
; 
32'd15786: dataIn1 = 32'd44
; 
32'd15787: dataIn1 = 32'd51
; 
32'd15788: dataIn1 = 32'd55
; 
32'd15789: dataIn1 = 32'd60
; 
32'd15790: dataIn1 = 32'd62
; 
32'd15791: dataIn1 = 32'd3
; 
32'd15792: dataIn1 = 32'd4
; 
32'd15793: dataIn1 = 32'd14
; 
32'd15794: dataIn1 = 32'd15
; 
32'd15795: dataIn1 = 32'd19
; 
32'd15796: dataIn1 = 32'd20
; 
32'd15797: dataIn1 = 32'd27
; 
32'd15798: dataIn1 = 32'd29
; 
32'd15799: dataIn1 = 32'd30
; 
32'd15800: dataIn1 = 32'd33
; 
32'd15801: dataIn1 = 32'd35
; 
32'd15802: dataIn1 = 32'd38
; 
32'd15803: dataIn1 = 32'd40
; 
32'd15804: dataIn1 = 32'd42
; 
32'd15805: dataIn1 = 32'd43
; 
32'd15806: dataIn1 = 32'd51
; 
32'd15807: dataIn1 = 32'd52
; 
32'd15808: dataIn1 = 32'd54
; 
32'd15809: dataIn1 = 32'd60
; 
32'd15810: dataIn1 = 32'd61
; 
32'd15811: dataIn1 = 32'd0
; 
32'd15812: dataIn1 = 32'd2
; 
32'd15813: dataIn1 = 32'd3
; 
32'd15814: dataIn1 = 32'd4
; 
32'd15815: dataIn1 = 32'd6
; 
32'd15816: dataIn1 = 32'd12
; 
32'd15817: dataIn1 = 32'd19
; 
32'd15818: dataIn1 = 32'd21
; 
32'd15819: dataIn1 = 32'd31
; 
32'd15820: dataIn1 = 32'd33
; 
32'd15821: dataIn1 = 32'd41
; 
32'd15822: dataIn1 = 32'd43
; 
32'd15823: dataIn1 = 32'd44
; 
32'd15824: dataIn1 = 32'd47
; 
32'd15825: dataIn1 = 32'd57
; 
32'd15826: dataIn1 = 32'd62
; 
32'd15827: dataIn1 = 32'd63
; 
32'd15828: dataIn1 = 32'd0
; 
32'd15829: dataIn1 = 32'd5
; 
32'd15830: dataIn1 = 32'd6
; 
32'd15831: dataIn1 = 32'd10
; 
32'd15832: dataIn1 = 32'd12
; 
32'd15833: dataIn1 = 32'd16
; 
32'd15834: dataIn1 = 32'd17
; 
32'd15835: dataIn1 = 32'd20
; 
32'd15836: dataIn1 = 32'd22
; 
32'd15837: dataIn1 = 32'd25
; 
32'd15838: dataIn1 = 32'd28
; 
32'd15839: dataIn1 = 32'd31
; 
32'd15840: dataIn1 = 32'd39
; 
32'd15841: dataIn1 = 32'd48
; 
32'd15842: dataIn1 = 32'd55
; 
32'd15843: dataIn1 = 32'd57
; 
32'd15844: dataIn1 = 32'd58
; 
32'd15845: dataIn1 = 32'd61
; 
32'd15846: dataIn1 = 32'd0
; 
32'd15847: dataIn1 = 32'd1
; 
32'd15848: dataIn1 = 32'd9
; 
32'd15849: dataIn1 = 32'd10
; 
32'd15850: dataIn1 = 32'd12
; 
32'd15851: dataIn1 = 32'd14
; 
32'd15852: dataIn1 = 32'd17
; 
32'd15853: dataIn1 = 32'd21
; 
32'd15854: dataIn1 = 32'd23
; 
32'd15855: dataIn1 = 32'd31
; 
32'd15856: dataIn1 = 32'd32
; 
32'd15857: dataIn1 = 32'd40
; 
32'd15858: dataIn1 = 32'd42
; 
32'd15859: dataIn1 = 32'd44
; 
32'd15860: dataIn1 = 32'd47
; 
32'd15861: dataIn1 = 32'd52
; 
32'd15862: dataIn1 = 32'd62
; 
32'd15863: dataIn1 = 32'd1
; 
32'd15864: dataIn1 = 32'd3
; 
32'd15865: dataIn1 = 32'd8
; 
32'd15866: dataIn1 = 32'd23
; 
32'd15867: dataIn1 = 32'd26
; 
32'd15868: dataIn1 = 32'd29
; 
32'd15869: dataIn1 = 32'd31
; 
32'd15870: dataIn1 = 32'd42
; 
32'd15871: dataIn1 = 32'd52
; 
32'd15872: dataIn1 = 32'd0
; 
32'd15873: dataIn1 = 32'd1
; 
32'd15874: dataIn1 = 32'd2
; 
32'd15875: dataIn1 = 32'd4
; 
32'd15876: dataIn1 = 32'd11
; 
32'd15877: dataIn1 = 32'd17
; 
32'd15878: dataIn1 = 32'd21
; 
32'd15879: dataIn1 = 32'd25
; 
32'd15880: dataIn1 = 32'd27
; 
32'd15881: dataIn1 = 32'd28
; 
32'd15882: dataIn1 = 32'd31
; 
32'd15883: dataIn1 = 32'd36
; 
32'd15884: dataIn1 = 32'd37
; 
32'd15885: dataIn1 = 32'd41
; 
32'd15886: dataIn1 = 32'd45
; 
32'd15887: dataIn1 = 32'd48
; 
32'd15888: dataIn1 = 32'd50
; 
32'd15889: dataIn1 = 32'd54
; 
32'd15890: dataIn1 = 32'd58
; 
32'd15891: dataIn1 = 32'd60
; 
32'd15892: dataIn1 = 32'd63
; 
32'd15893: dataIn1 = 32'd1
; 
32'd15894: dataIn1 = 32'd4
; 
32'd15895: dataIn1 = 32'd7
; 
32'd15896: dataIn1 = 32'd11
; 
32'd15897: dataIn1 = 32'd15
; 
32'd15898: dataIn1 = 32'd16
; 
32'd15899: dataIn1 = 32'd23
; 
32'd15900: dataIn1 = 32'd32
; 
32'd15901: dataIn1 = 32'd33
; 
32'd15902: dataIn1 = 32'd37
; 
32'd15903: dataIn1 = 32'd44
; 
32'd15904: dataIn1 = 32'd45
; 
32'd15905: dataIn1 = 32'd46
; 
32'd15906: dataIn1 = 32'd49
; 
32'd15907: dataIn1 = 32'd53
; 
32'd15908: dataIn1 = 32'd56
; 
32'd15909: dataIn1 = 32'd57
; 
32'd15910: dataIn1 = 32'd63
; 
32'd15911: dataIn1 = 32'd6
; 
32'd15912: dataIn1 = 32'd8
; 
32'd15913: dataIn1 = 32'd13
; 
32'd15914: dataIn1 = 32'd16
; 
32'd15915: dataIn1 = 32'd18
; 
32'd15916: dataIn1 = 32'd24
; 
32'd15917: dataIn1 = 32'd26
; 
32'd15918: dataIn1 = 32'd27
; 
32'd15919: dataIn1 = 32'd33
; 
32'd15920: dataIn1 = 32'd37
; 
32'd15921: dataIn1 = 32'd38
; 
32'd15922: dataIn1 = 32'd41
; 
32'd15923: dataIn1 = 32'd44
; 
32'd15924: dataIn1 = 32'd45
; 
32'd15925: dataIn1 = 32'd53
; 
32'd15926: dataIn1 = 32'd56
; 
32'd15927: dataIn1 = 32'd58
; 
32'd15928: dataIn1 = 32'd60
; 
32'd15929: dataIn1 = 32'd61
; 
32'd15930: dataIn1 = 32'd63
; 
32'd15931: dataIn1 = 32'd3
; 
32'd15932: dataIn1 = 32'd4
; 
32'd15933: dataIn1 = 32'd8
; 
32'd15934: dataIn1 = 32'd9
; 
32'd15935: dataIn1 = 32'd16
; 
32'd15936: dataIn1 = 32'd20
; 
32'd15937: dataIn1 = 32'd22
; 
32'd15938: dataIn1 = 32'd27
; 
32'd15939: dataIn1 = 32'd30
; 
32'd15940: dataIn1 = 32'd31
; 
32'd15941: dataIn1 = 32'd33
; 
32'd15942: dataIn1 = 32'd35
; 
32'd15943: dataIn1 = 32'd39
; 
32'd15944: dataIn1 = 32'd40
; 
32'd15945: dataIn1 = 32'd41
; 
32'd15946: dataIn1 = 32'd46
; 
32'd15947: dataIn1 = 32'd47
; 
32'd15948: dataIn1 = 32'd49
; 
32'd15949: dataIn1 = 32'd51
; 
32'd15950: dataIn1 = 32'd56
; 
32'd15951: dataIn1 = 32'd60
; 
32'd15952: dataIn1 = 32'd11
; 
32'd15953: dataIn1 = 32'd12
; 
32'd15954: dataIn1 = 32'd16
; 
32'd15955: dataIn1 = 32'd21
; 
32'd15956: dataIn1 = 32'd24
; 
32'd15957: dataIn1 = 32'd26
; 
32'd15958: dataIn1 = 32'd30
; 
32'd15959: dataIn1 = 32'd32
; 
32'd15960: dataIn1 = 32'd33
; 
32'd15961: dataIn1 = 32'd40
; 
32'd15962: dataIn1 = 32'd47
; 
32'd15963: dataIn1 = 32'd50
; 
32'd15964: dataIn1 = 32'd51
; 
32'd15965: dataIn1 = 32'd54
; 
32'd15966: dataIn1 = 32'd56
; 
32'd15967: dataIn1 = 32'd61
; 
32'd15968: dataIn1 = 32'd0
; 
32'd15969: dataIn1 = 32'd4
; 
32'd15970: dataIn1 = 32'd5
; 
32'd15971: dataIn1 = 32'd6
; 
32'd15972: dataIn1 = 32'd10
; 
32'd15973: dataIn1 = 32'd12
; 
32'd15974: dataIn1 = 32'd17
; 
32'd15975: dataIn1 = 32'd26
; 
32'd15976: dataIn1 = 32'd27
; 
32'd15977: dataIn1 = 32'd28
; 
32'd15978: dataIn1 = 32'd29
; 
32'd15979: dataIn1 = 32'd30
; 
32'd15980: dataIn1 = 32'd37
; 
32'd15981: dataIn1 = 32'd39
; 
32'd15982: dataIn1 = 32'd41
; 
32'd15983: dataIn1 = 32'd42
; 
32'd15984: dataIn1 = 32'd51
; 
32'd15985: dataIn1 = 32'd52
; 
32'd15986: dataIn1 = 32'd54
; 
32'd15987: dataIn1 = 32'd60
; 
32'd15988: dataIn1 = 32'd62
; 
32'd15989: dataIn1 = 32'd3
; 
32'd15990: dataIn1 = 32'd5
; 
32'd15991: dataIn1 = 32'd14
; 
32'd15992: dataIn1 = 32'd16
; 
32'd15993: dataIn1 = 32'd18
; 
32'd15994: dataIn1 = 32'd20
; 
32'd15995: dataIn1 = 32'd21
; 
32'd15996: dataIn1 = 32'd24
; 
32'd15997: dataIn1 = 32'd28
; 
32'd15998: dataIn1 = 32'd30
; 
32'd15999: dataIn1 = 32'd46
; 
32'd16000: dataIn1 = 32'd47
; 
32'd16001: dataIn1 = 32'd49
; 
32'd16002: dataIn1 = 32'd51
; 
32'd16003: dataIn1 = 32'd55
; 
32'd16004: dataIn1 = 32'd56
; 
32'd16005: dataIn1 = 32'd57
; 
32'd16006: dataIn1 = 32'd58
; 
32'd16007: dataIn1 = 32'd62
; 
32'd16008: dataIn1 = 32'd63
; 
32'd16009: dataIn1 = 32'd0
; 
32'd16010: dataIn1 = 32'd1
; 
32'd16011: dataIn1 = 32'd5
; 
32'd16012: dataIn1 = 32'd6
; 
32'd16013: dataIn1 = 32'd8
; 
32'd16014: dataIn1 = 32'd11
; 
32'd16015: dataIn1 = 32'd20
; 
32'd16016: dataIn1 = 32'd21
; 
32'd16017: dataIn1 = 32'd22
; 
32'd16018: dataIn1 = 32'd24
; 
32'd16019: dataIn1 = 32'd32
; 
32'd16020: dataIn1 = 32'd33
; 
32'd16021: dataIn1 = 32'd34
; 
32'd16022: dataIn1 = 32'd35
; 
32'd16023: dataIn1 = 32'd38
; 
32'd16024: dataIn1 = 32'd40
; 
32'd16025: dataIn1 = 32'd44
; 
32'd16026: dataIn1 = 32'd45
; 
32'd16027: dataIn1 = 32'd46
; 
32'd16028: dataIn1 = 32'd49
; 
32'd16029: dataIn1 = 32'd53
; 
32'd16030: dataIn1 = 32'd55
; 
32'd16031: dataIn1 = 32'd59
; 
32'd16032: dataIn1 = 32'd63
; 
32'd16033: dataIn1 = 32'd3
; 
32'd16034: dataIn1 = 32'd7
; 
32'd16035: dataIn1 = 32'd15
; 
32'd16036: dataIn1 = 32'd16
; 
32'd16037: dataIn1 = 32'd20
; 
32'd16038: dataIn1 = 32'd21
; 
32'd16039: dataIn1 = 32'd22
; 
32'd16040: dataIn1 = 32'd23
; 
32'd16041: dataIn1 = 32'd24
; 
32'd16042: dataIn1 = 32'd25
; 
32'd16043: dataIn1 = 32'd29
; 
32'd16044: dataIn1 = 32'd31
; 
32'd16045: dataIn1 = 32'd38
; 
32'd16046: dataIn1 = 32'd39
; 
32'd16047: dataIn1 = 32'd41
; 
32'd16048: dataIn1 = 32'd43
; 
32'd16049: dataIn1 = 32'd51
; 
32'd16050: dataIn1 = 32'd52
; 
32'd16051: dataIn1 = 32'd53
; 
32'd16052: dataIn1 = 32'd58
; 
32'd16053: dataIn1 = 32'd59
; 
32'd16054: dataIn1 = 32'd0
; 
32'd16055: dataIn1 = 32'd4
; 
32'd16056: dataIn1 = 32'd5
; 
32'd16057: dataIn1 = 32'd7
; 
32'd16058: dataIn1 = 32'd9
; 
32'd16059: dataIn1 = 32'd11
; 
32'd16060: dataIn1 = 32'd12
; 
32'd16061: dataIn1 = 32'd14
; 
32'd16062: dataIn1 = 32'd17
; 
32'd16063: dataIn1 = 32'd18
; 
32'd16064: dataIn1 = 32'd23
; 
32'd16065: dataIn1 = 32'd30
; 
32'd16066: dataIn1 = 32'd31
; 
32'd16067: dataIn1 = 32'd34
; 
32'd16068: dataIn1 = 32'd35
; 
32'd16069: dataIn1 = 32'd42
; 
32'd16070: dataIn1 = 32'd44
; 
32'd16071: dataIn1 = 32'd52
; 
32'd16072: dataIn1 = 32'd55
; 
32'd16073: dataIn1 = 32'd56
; 
32'd16074: dataIn1 = 32'd59
; 
32'd16075: dataIn1 = 32'd63
; 
32'd16076: dataIn1 = 32'd1
; 
32'd16077: dataIn1 = 32'd8
; 
32'd16078: dataIn1 = 32'd10
; 
32'd16079: dataIn1 = 32'd21
; 
32'd16080: dataIn1 = 32'd23
; 
32'd16081: dataIn1 = 32'd34
; 
32'd16082: dataIn1 = 32'd35
; 
32'd16083: dataIn1 = 32'd36
; 
32'd16084: dataIn1 = 32'd37
; 
32'd16085: dataIn1 = 32'd41
; 
32'd16086: dataIn1 = 32'd43
; 
32'd16087: dataIn1 = 32'd47
; 
32'd16088: dataIn1 = 32'd51
; 
32'd16089: dataIn1 = 32'd52
; 
32'd16090: dataIn1 = 32'd53
; 
32'd16091: dataIn1 = 32'd4
; 
32'd16092: dataIn1 = 32'd5
; 
32'd16093: dataIn1 = 32'd9
; 
32'd16094: dataIn1 = 32'd12
; 
32'd16095: dataIn1 = 32'd17
; 
32'd16096: dataIn1 = 32'd20
; 
32'd16097: dataIn1 = 32'd21
; 
32'd16098: dataIn1 = 32'd24
; 
32'd16099: dataIn1 = 32'd25
; 
32'd16100: dataIn1 = 32'd35
; 
32'd16101: dataIn1 = 32'd39
; 
32'd16102: dataIn1 = 32'd44
; 
32'd16103: dataIn1 = 32'd55
; 
32'd16104: dataIn1 = 32'd56
; 
32'd16105: dataIn1 = 32'd57
; 
32'd16106: dataIn1 = 32'd58
; 
32'd16107: dataIn1 = 32'd62
; 
32'd16108: dataIn1 = 32'd63
; 
32'd16109: dataIn1 = 32'd0
; 
32'd16110: dataIn1 = 32'd2
; 
32'd16111: dataIn1 = 32'd3
; 
32'd16112: dataIn1 = 32'd6
; 
32'd16113: dataIn1 = 32'd7
; 
32'd16114: dataIn1 = 32'd13
; 
32'd16115: dataIn1 = 32'd18
; 
32'd16116: dataIn1 = 32'd19
; 
32'd16117: dataIn1 = 32'd21
; 
32'd16118: dataIn1 = 32'd25
; 
32'd16119: dataIn1 = 32'd29
; 
32'd16120: dataIn1 = 32'd30
; 
32'd16121: dataIn1 = 32'd35
; 
32'd16122: dataIn1 = 32'd36
; 
32'd16123: dataIn1 = 32'd37
; 
32'd16124: dataIn1 = 32'd38
; 
32'd16125: dataIn1 = 32'd39
; 
32'd16126: dataIn1 = 32'd42
; 
32'd16127: dataIn1 = 32'd46
; 
32'd16128: dataIn1 = 32'd47
; 
32'd16129: dataIn1 = 32'd49
; 
32'd16130: dataIn1 = 32'd50
; 
32'd16131: dataIn1 = 32'd51
; 
32'd16132: dataIn1 = 32'd53
; 
32'd16133: dataIn1 = 32'd56
; 
32'd16134: dataIn1 = 32'd60
; 
32'd16135: dataIn1 = 32'd62
; 
32'd16136: dataIn1 = 32'd63
; 
32'd16137: dataIn1 = 32'd1
; 
32'd16138: dataIn1 = 32'd2
; 
32'd16139: dataIn1 = 32'd10
; 
32'd16140: dataIn1 = 32'd12
; 
32'd16141: dataIn1 = 32'd13
; 
32'd16142: dataIn1 = 32'd17
; 
32'd16143: dataIn1 = 32'd18
; 
32'd16144: dataIn1 = 32'd19
; 
32'd16145: dataIn1 = 32'd25
; 
32'd16146: dataIn1 = 32'd32
; 
32'd16147: dataIn1 = 32'd36
; 
32'd16148: dataIn1 = 32'd43
; 
32'd16149: dataIn1 = 32'd44
; 
32'd16150: dataIn1 = 32'd47
; 
32'd16151: dataIn1 = 32'd50
; 
32'd16152: dataIn1 = 32'd51
; 
32'd16153: dataIn1 = 32'd1
; 
32'd16154: dataIn1 = 32'd2
; 
32'd16155: dataIn1 = 32'd5
; 
32'd16156: dataIn1 = 32'd6
; 
32'd16157: dataIn1 = 32'd7
; 
32'd16158: dataIn1 = 32'd8
; 
32'd16159: dataIn1 = 32'd10
; 
32'd16160: dataIn1 = 32'd12
; 
32'd16161: dataIn1 = 32'd14
; 
32'd16162: dataIn1 = 32'd18
; 
32'd16163: dataIn1 = 32'd23
; 
32'd16164: dataIn1 = 32'd28
; 
32'd16165: dataIn1 = 32'd30
; 
32'd16166: dataIn1 = 32'd32
; 
32'd16167: dataIn1 = 32'd36
; 
32'd16168: dataIn1 = 32'd40
; 
32'd16169: dataIn1 = 32'd44
; 
32'd16170: dataIn1 = 32'd47
; 
32'd16171: dataIn1 = 32'd56
; 
32'd16172: dataIn1 = 32'd61
; 
32'd16173: dataIn1 = 32'd2
; 
32'd16174: dataIn1 = 32'd3
; 
32'd16175: dataIn1 = 32'd5
; 
32'd16176: dataIn1 = 32'd7
; 
32'd16177: dataIn1 = 32'd10
; 
32'd16178: dataIn1 = 32'd15
; 
32'd16179: dataIn1 = 32'd17
; 
32'd16180: dataIn1 = 32'd18
; 
32'd16181: dataIn1 = 32'd29
; 
32'd16182: dataIn1 = 32'd34
; 
32'd16183: dataIn1 = 32'd35
; 
32'd16184: dataIn1 = 32'd36
; 
32'd16185: dataIn1 = 32'd40
; 
32'd16186: dataIn1 = 32'd42
; 
32'd16187: dataIn1 = 32'd43
; 
32'd16188: dataIn1 = 32'd44
; 
32'd16189: dataIn1 = 32'd51
; 
32'd16190: dataIn1 = 32'd55
; 
32'd16191: dataIn1 = 32'd4
; 
32'd16192: dataIn1 = 32'd11
; 
32'd16193: dataIn1 = 32'd14
; 
32'd16194: dataIn1 = 32'd15
; 
32'd16195: dataIn1 = 32'd26
; 
32'd16196: dataIn1 = 32'd27
; 
32'd16197: dataIn1 = 32'd28
; 
32'd16198: dataIn1 = 32'd30
; 
32'd16199: dataIn1 = 32'd36
; 
32'd16200: dataIn1 = 32'd41
; 
32'd16201: dataIn1 = 32'd42
; 
32'd16202: dataIn1 = 32'd46
; 
32'd16203: dataIn1 = 32'd48
; 
32'd16204: dataIn1 = 32'd54
; 
32'd16205: dataIn1 = 32'd58
; 
32'd16206: dataIn1 = 32'd2
; 
32'd16207: dataIn1 = 32'd6
; 
32'd16208: dataIn1 = 32'd7
; 
32'd16209: dataIn1 = 32'd9
; 
32'd16210: dataIn1 = 32'd13
; 
32'd16211: dataIn1 = 32'd14
; 
32'd16212: dataIn1 = 32'd15
; 
32'd16213: dataIn1 = 32'd19
; 
32'd16214: dataIn1 = 32'd22
; 
32'd16215: dataIn1 = 32'd24
; 
32'd16216: dataIn1 = 32'd27
; 
32'd16217: dataIn1 = 32'd35
; 
32'd16218: dataIn1 = 32'd37
; 
32'd16219: dataIn1 = 32'd44
; 
32'd16220: dataIn1 = 32'd50
; 
32'd16221: dataIn1 = 32'd51
; 
32'd16222: dataIn1 = 32'd54
; 
32'd16223: dataIn1 = 32'd63
; 
32'd16224: dataIn1 = 32'd3
; 
32'd16225: dataIn1 = 32'd5
; 
32'd16226: dataIn1 = 32'd9
; 
32'd16227: dataIn1 = 32'd11
; 
32'd16228: dataIn1 = 32'd14
; 
32'd16229: dataIn1 = 32'd15
; 
32'd16230: dataIn1 = 32'd24
; 
32'd16231: dataIn1 = 32'd26
; 
32'd16232: dataIn1 = 32'd32
; 
32'd16233: dataIn1 = 32'd33
; 
32'd16234: dataIn1 = 32'd37
; 
32'd16235: dataIn1 = 32'd38
; 
32'd16236: dataIn1 = 32'd41
; 
32'd16237: dataIn1 = 32'd43
; 
32'd16238: dataIn1 = 32'd46
; 
32'd16239: dataIn1 = 32'd50
; 
32'd16240: dataIn1 = 32'd54
; 
32'd16241: dataIn1 = 32'd55
; 
32'd16242: dataIn1 = 32'd60
; 
32'd16243: dataIn1 = 32'd0
; 
32'd16244: dataIn1 = 32'd7
; 
32'd16245: dataIn1 = 32'd12
; 
32'd16246: dataIn1 = 32'd19
; 
32'd16247: dataIn1 = 32'd26
; 
32'd16248: dataIn1 = 32'd31
; 
32'd16249: dataIn1 = 32'd34
; 
32'd16250: dataIn1 = 32'd37
; 
32'd16251: dataIn1 = 32'd38
; 
32'd16252: dataIn1 = 32'd43
; 
32'd16253: dataIn1 = 32'd49
; 
32'd16254: dataIn1 = 32'd52
; 
32'd16255: dataIn1 = 32'd55
; 
32'd16256: dataIn1 = 32'd60
; 
32'd16257: dataIn1 = 32'd63
; 
32'd16258: dataIn1 = 32'd1
; 
32'd16259: dataIn1 = 32'd2
; 
32'd16260: dataIn1 = 32'd3
; 
32'd16261: dataIn1 = 32'd4
; 
32'd16262: dataIn1 = 32'd6
; 
32'd16263: dataIn1 = 32'd10
; 
32'd16264: dataIn1 = 32'd11
; 
32'd16265: dataIn1 = 32'd26
; 
32'd16266: dataIn1 = 32'd28
; 
32'd16267: dataIn1 = 32'd29
; 
32'd16268: dataIn1 = 32'd30
; 
32'd16269: dataIn1 = 32'd32
; 
32'd16270: dataIn1 = 32'd34
; 
32'd16271: dataIn1 = 32'd37
; 
32'd16272: dataIn1 = 32'd39
; 
32'd16273: dataIn1 = 32'd42
; 
32'd16274: dataIn1 = 32'd45
; 
32'd16275: dataIn1 = 32'd56
; 
32'd16276: dataIn1 = 32'd57
; 
32'd16277: dataIn1 = 32'd59
; 
32'd16278: dataIn1 = 32'd4
; 
32'd16279: dataIn1 = 32'd11
; 
32'd16280: dataIn1 = 32'd16
; 
32'd16281: dataIn1 = 32'd22
; 
32'd16282: dataIn1 = 32'd24
; 
32'd16283: dataIn1 = 32'd28
; 
32'd16284: dataIn1 = 32'd31
; 
32'd16285: dataIn1 = 32'd32
; 
32'd16286: dataIn1 = 32'd35
; 
32'd16287: dataIn1 = 32'd36
; 
32'd16288: dataIn1 = 32'd38
; 
32'd16289: dataIn1 = 32'd56
; 
32'd16290: dataIn1 = 32'd61
; 
32'd16291: dataIn1 = 32'd63
; 
32'd16292: dataIn1 = 32'd0
; 
32'd16293: dataIn1 = 32'd6
; 
32'd16294: dataIn1 = 32'd8
; 
32'd16295: dataIn1 = 32'd18
; 
32'd16296: dataIn1 = 32'd26
; 
32'd16297: dataIn1 = 32'd28
; 
32'd16298: dataIn1 = 32'd32
; 
32'd16299: dataIn1 = 32'd34
; 
32'd16300: dataIn1 = 32'd35
; 
32'd16301: dataIn1 = 32'd37
; 
32'd16302: dataIn1 = 32'd38
; 
32'd16303: dataIn1 = 32'd41
; 
32'd16304: dataIn1 = 32'd42
; 
32'd16305: dataIn1 = 32'd45
; 
32'd16306: dataIn1 = 32'd50
; 
32'd16307: dataIn1 = 32'd55
; 
32'd16308: dataIn1 = 32'd57
; 
32'd16309: dataIn1 = 32'd61
; 
32'd16310: dataIn1 = 32'd5
; 
32'd16311: dataIn1 = 32'd15
; 
32'd16312: dataIn1 = 32'd21
; 
32'd16313: dataIn1 = 32'd22
; 
32'd16314: dataIn1 = 32'd23
; 
32'd16315: dataIn1 = 32'd28
; 
32'd16316: dataIn1 = 32'd30
; 
32'd16317: dataIn1 = 32'd32
; 
32'd16318: dataIn1 = 32'd33
; 
32'd16319: dataIn1 = 32'd39
; 
32'd16320: dataIn1 = 32'd41
; 
32'd16321: dataIn1 = 32'd44
; 
32'd16322: dataIn1 = 32'd50
; 
32'd16323: dataIn1 = 32'd52
; 
32'd16324: dataIn1 = 32'd56
; 
32'd16325: dataIn1 = 32'd59
; 
32'd16326: dataIn1 = 32'd62
; 
32'd16327: dataIn1 = 32'd2
; 
32'd16328: dataIn1 = 32'd4
; 
32'd16329: dataIn1 = 32'd10
; 
32'd16330: dataIn1 = 32'd11
; 
32'd16331: dataIn1 = 32'd16
; 
32'd16332: dataIn1 = 32'd22
; 
32'd16333: dataIn1 = 32'd28
; 
32'd16334: dataIn1 = 32'd30
; 
32'd16335: dataIn1 = 32'd36
; 
32'd16336: dataIn1 = 32'd43
; 
32'd16337: dataIn1 = 32'd44
; 
32'd16338: dataIn1 = 32'd45
; 
32'd16339: dataIn1 = 32'd50
; 
32'd16340: dataIn1 = 32'd51
; 
32'd16341: dataIn1 = 32'd52
; 
32'd16342: dataIn1 = 32'd53
; 
32'd16343: dataIn1 = 32'd57
; 
32'd16344: dataIn1 = 32'd58
; 
32'd16345: dataIn1 = 32'd59
; 
32'd16346: dataIn1 = 32'd60
; 
32'd16347: dataIn1 = 32'd62
; 
32'd16348: dataIn1 = 32'd4
; 
32'd16349: dataIn1 = 32'd7
; 
32'd16350: dataIn1 = 32'd10
; 
32'd16351: dataIn1 = 32'd14
; 
32'd16352: dataIn1 = 32'd15
; 
32'd16353: dataIn1 = 32'd16
; 
32'd16354: dataIn1 = 32'd17
; 
32'd16355: dataIn1 = 32'd20
; 
32'd16356: dataIn1 = 32'd34
; 
32'd16357: dataIn1 = 32'd39
; 
32'd16358: dataIn1 = 32'd43
; 
32'd16359: dataIn1 = 32'd47
; 
32'd16360: dataIn1 = 32'd54
; 
32'd16361: dataIn1 = 32'd57
; 
32'd16362: dataIn1 = 32'd0
; 
32'd16363: dataIn1 = 32'd1
; 
32'd16364: dataIn1 = 32'd4
; 
32'd16365: dataIn1 = 32'd9
; 
32'd16366: dataIn1 = 32'd11
; 
32'd16367: dataIn1 = 32'd16
; 
32'd16368: dataIn1 = 32'd21
; 
32'd16369: dataIn1 = 32'd30
; 
32'd16370: dataIn1 = 32'd36
; 
32'd16371: dataIn1 = 32'd38
; 
32'd16372: dataIn1 = 32'd40
; 
32'd16373: dataIn1 = 32'd44
; 
32'd16374: dataIn1 = 32'd47
; 
32'd16375: dataIn1 = 32'd50
; 
32'd16376: dataIn1 = 32'd53
; 
32'd16377: dataIn1 = 32'd59
; 
32'd16378: dataIn1 = 32'd62
; 
32'd16379: dataIn1 = 32'd1
; 
32'd16380: dataIn1 = 32'd4
; 
32'd16381: dataIn1 = 32'd6
; 
32'd16382: dataIn1 = 32'd18
; 
32'd16383: dataIn1 = 32'd26
; 
32'd16384: dataIn1 = 32'd30
; 
32'd16385: dataIn1 = 32'd31
; 
32'd16386: dataIn1 = 32'd33
; 
32'd16387: dataIn1 = 32'd34
; 
32'd16388: dataIn1 = 32'd39
; 
32'd16389: dataIn1 = 32'd41
; 
32'd16390: dataIn1 = 32'd44
; 
32'd16391: dataIn1 = 32'd45
; 
32'd16392: dataIn1 = 32'd49
; 
32'd16393: dataIn1 = 32'd51
; 
32'd16394: dataIn1 = 32'd55
; 
32'd16395: dataIn1 = 32'd2
; 
32'd16396: dataIn1 = 32'd3
; 
32'd16397: dataIn1 = 32'd4
; 
32'd16398: dataIn1 = 32'd6
; 
32'd16399: dataIn1 = 32'd7
; 
32'd16400: dataIn1 = 32'd8
; 
32'd16401: dataIn1 = 32'd11
; 
32'd16402: dataIn1 = 32'd12
; 
32'd16403: dataIn1 = 32'd18
; 
32'd16404: dataIn1 = 32'd24
; 
32'd16405: dataIn1 = 32'd30
; 
32'd16406: dataIn1 = 32'd36
; 
32'd16407: dataIn1 = 32'd40
; 
32'd16408: dataIn1 = 32'd44
; 
32'd16409: dataIn1 = 32'd49
; 
32'd16410: dataIn1 = 32'd53
; 
32'd16411: dataIn1 = 32'd54
; 
32'd16412: dataIn1 = 32'd57
; 
32'd16413: dataIn1 = 32'd61
; 
32'd16414: dataIn1 = 32'd62
; 
32'd16415: dataIn1 = 32'd63
; 
32'd16416: dataIn1 = 32'd2
; 
32'd16417: dataIn1 = 32'd3
; 
32'd16418: dataIn1 = 32'd5
; 
32'd16419: dataIn1 = 32'd6
; 
32'd16420: dataIn1 = 32'd7
; 
32'd16421: dataIn1 = 32'd23
; 
32'd16422: dataIn1 = 32'd26
; 
32'd16423: dataIn1 = 32'd30
; 
32'd16424: dataIn1 = 32'd32
; 
32'd16425: dataIn1 = 32'd35
; 
32'd16426: dataIn1 = 32'd39
; 
32'd16427: dataIn1 = 32'd41
; 
32'd16428: dataIn1 = 32'd44
; 
32'd16429: dataIn1 = 32'd56
; 
32'd16430: dataIn1 = 32'd63
; 
32'd16431: dataIn1 = 32'd0
; 
32'd16432: dataIn1 = 32'd3
; 
32'd16433: dataIn1 = 32'd4
; 
32'd16434: dataIn1 = 32'd7
; 
32'd16435: dataIn1 = 32'd16
; 
32'd16436: dataIn1 = 32'd18
; 
32'd16437: dataIn1 = 32'd22
; 
32'd16438: dataIn1 = 32'd23
; 
32'd16439: dataIn1 = 32'd24
; 
32'd16440: dataIn1 = 32'd25
; 
32'd16441: dataIn1 = 32'd33
; 
32'd16442: dataIn1 = 32'd34
; 
32'd16443: dataIn1 = 32'd35
; 
32'd16444: dataIn1 = 32'd36
; 
32'd16445: dataIn1 = 32'd38
; 
32'd16446: dataIn1 = 32'd40
; 
32'd16447: dataIn1 = 32'd44
; 
32'd16448: dataIn1 = 32'd45
; 
32'd16449: dataIn1 = 32'd46
; 
32'd16450: dataIn1 = 32'd53
; 
32'd16451: dataIn1 = 32'd56
; 
32'd16452: dataIn1 = 32'd61
; 
32'd16453: dataIn1 = 32'd62
; 
32'd16454: dataIn1 = 32'd1
; 
32'd16455: dataIn1 = 32'd2
; 
32'd16456: dataIn1 = 32'd4
; 
32'd16457: dataIn1 = 32'd7
; 
32'd16458: dataIn1 = 32'd11
; 
32'd16459: dataIn1 = 32'd12
; 
32'd16460: dataIn1 = 32'd13
; 
32'd16461: dataIn1 = 32'd21
; 
32'd16462: dataIn1 = 32'd31
; 
32'd16463: dataIn1 = 32'd34
; 
32'd16464: dataIn1 = 32'd36
; 
32'd16465: dataIn1 = 32'd38
; 
32'd16466: dataIn1 = 32'd41
; 
32'd16467: dataIn1 = 32'd48
; 
32'd16468: dataIn1 = 32'd50
; 
32'd16469: dataIn1 = 32'd53
; 
32'd16470: dataIn1 = 32'd59
; 
32'd16471: dataIn1 = 32'd60
; 
32'd16472: dataIn1 = 32'd1
; 
32'd16473: dataIn1 = 32'd4
; 
32'd16474: dataIn1 = 32'd9
; 
32'd16475: dataIn1 = 32'd11
; 
32'd16476: dataIn1 = 32'd17
; 
32'd16477: dataIn1 = 32'd18
; 
32'd16478: dataIn1 = 32'd20
; 
32'd16479: dataIn1 = 32'd21
; 
32'd16480: dataIn1 = 32'd22
; 
32'd16481: dataIn1 = 32'd24
; 
32'd16482: dataIn1 = 32'd25
; 
32'd16483: dataIn1 = 32'd27
; 
32'd16484: dataIn1 = 32'd32
; 
32'd16485: dataIn1 = 32'd34
; 
32'd16486: dataIn1 = 32'd35
; 
32'd16487: dataIn1 = 32'd43
; 
32'd16488: dataIn1 = 32'd45
; 
32'd16489: dataIn1 = 32'd48
; 
32'd16490: dataIn1 = 32'd49
; 
32'd16491: dataIn1 = 32'd50
; 
32'd16492: dataIn1 = 32'd56
; 
32'd16493: dataIn1 = 32'd58
; 
32'd16494: dataIn1 = 32'd62
; 
32'd16495: dataIn1 = 32'd1
; 
32'd16496: dataIn1 = 32'd2
; 
32'd16497: dataIn1 = 32'd10
; 
32'd16498: dataIn1 = 32'd15
; 
32'd16499: dataIn1 = 32'd16
; 
32'd16500: dataIn1 = 32'd17
; 
32'd16501: dataIn1 = 32'd18
; 
32'd16502: dataIn1 = 32'd22
; 
32'd16503: dataIn1 = 32'd26
; 
32'd16504: dataIn1 = 32'd28
; 
32'd16505: dataIn1 = 32'd29
; 
32'd16506: dataIn1 = 32'd37
; 
32'd16507: dataIn1 = 32'd51
; 
32'd16508: dataIn1 = 32'd54
; 
32'd16509: dataIn1 = 32'd61
; 
32'd16510: dataIn1 = 32'd7
; 
32'd16511: dataIn1 = 32'd8
; 
32'd16512: dataIn1 = 32'd11
; 
32'd16513: dataIn1 = 32'd13
; 
32'd16514: dataIn1 = 32'd16
; 
32'd16515: dataIn1 = 32'd17
; 
32'd16516: dataIn1 = 32'd22
; 
32'd16517: dataIn1 = 32'd23
; 
32'd16518: dataIn1 = 32'd24
; 
32'd16519: dataIn1 = 32'd26
; 
32'd16520: dataIn1 = 32'd27
; 
32'd16521: dataIn1 = 32'd28
; 
32'd16522: dataIn1 = 32'd31
; 
32'd16523: dataIn1 = 32'd34
; 
32'd16524: dataIn1 = 32'd39
; 
32'd16525: dataIn1 = 32'd41
; 
32'd16526: dataIn1 = 32'd42
; 
32'd16527: dataIn1 = 32'd46
; 
32'd16528: dataIn1 = 32'd49
; 
32'd16529: dataIn1 = 32'd50
; 
32'd16530: dataIn1 = 32'd54
; 
32'd16531: dataIn1 = 32'd55
; 
32'd16532: dataIn1 = 32'd58
; 
32'd16533: dataIn1 = 32'd59
; 
32'd16534: dataIn1 = 32'd61
; 
32'd16535: dataIn1 = 32'd1
; 
32'd16536: dataIn1 = 32'd6
; 
32'd16537: dataIn1 = 32'd11
; 
32'd16538: dataIn1 = 32'd12
; 
32'd16539: dataIn1 = 32'd17
; 
32'd16540: dataIn1 = 32'd21
; 
32'd16541: dataIn1 = 32'd23
; 
32'd16542: dataIn1 = 32'd24
; 
32'd16543: dataIn1 = 32'd31
; 
32'd16544: dataIn1 = 32'd34
; 
32'd16545: dataIn1 = 32'd37
; 
32'd16546: dataIn1 = 32'd38
; 
32'd16547: dataIn1 = 32'd40
; 
32'd16548: dataIn1 = 32'd45
; 
32'd16549: dataIn1 = 32'd46
; 
32'd16550: dataIn1 = 32'd48
; 
32'd16551: dataIn1 = 32'd49
; 
32'd16552: dataIn1 = 32'd50
; 
32'd16553: dataIn1 = 32'd62
; 
32'd16554: dataIn1 = 32'd6
; 
32'd16555: dataIn1 = 32'd17
; 
32'd16556: dataIn1 = 32'd18
; 
32'd16557: dataIn1 = 32'd20
; 
32'd16558: dataIn1 = 32'd23
; 
32'd16559: dataIn1 = 32'd24
; 
32'd16560: dataIn1 = 32'd26
; 
32'd16561: dataIn1 = 32'd29
; 
32'd16562: dataIn1 = 32'd31
; 
32'd16563: dataIn1 = 32'd34
; 
32'd16564: dataIn1 = 32'd42
; 
32'd16565: dataIn1 = 32'd44
; 
32'd16566: dataIn1 = 32'd46
; 
32'd16567: dataIn1 = 32'd47
; 
32'd16568: dataIn1 = 32'd52
; 
32'd16569: dataIn1 = 32'd61
; 
32'd16570: dataIn1 = 32'd62
; 
32'd16571: dataIn1 = 32'd2
; 
32'd16572: dataIn1 = 32'd8
; 
32'd16573: dataIn1 = 32'd10
; 
32'd16574: dataIn1 = 32'd11
; 
32'd16575: dataIn1 = 32'd12
; 
32'd16576: dataIn1 = 32'd13
; 
32'd16577: dataIn1 = 32'd18
; 
32'd16578: dataIn1 = 32'd22
; 
32'd16579: dataIn1 = 32'd24
; 
32'd16580: dataIn1 = 32'd27
; 
32'd16581: dataIn1 = 32'd29
; 
32'd16582: dataIn1 = 32'd32
; 
32'd16583: dataIn1 = 32'd35
; 
32'd16584: dataIn1 = 32'd39
; 
32'd16585: dataIn1 = 32'd45
; 
32'd16586: dataIn1 = 32'd50
; 
32'd16587: dataIn1 = 32'd60
; 
32'd16588: dataIn1 = 32'd61
; 
32'd16589: dataIn1 = 32'd3
; 
32'd16590: dataIn1 = 32'd9
; 
32'd16591: dataIn1 = 32'd15
; 
32'd16592: dataIn1 = 32'd17
; 
32'd16593: dataIn1 = 32'd19
; 
32'd16594: dataIn1 = 32'd26
; 
32'd16595: dataIn1 = 32'd35
; 
32'd16596: dataIn1 = 32'd39
; 
32'd16597: dataIn1 = 32'd41
; 
32'd16598: dataIn1 = 32'd45
; 
32'd16599: dataIn1 = 32'd47
; 
32'd16600: dataIn1 = 32'd53
; 
32'd16601: dataIn1 = 32'd5
; 
32'd16602: dataIn1 = 32'd7
; 
32'd16603: dataIn1 = 32'd9
; 
32'd16604: dataIn1 = 32'd14
; 
32'd16605: dataIn1 = 32'd16
; 
32'd16606: dataIn1 = 32'd19
; 
32'd16607: dataIn1 = 32'd21
; 
32'd16608: dataIn1 = 32'd22
; 
32'd16609: dataIn1 = 32'd24
; 
32'd16610: dataIn1 = 32'd30
; 
32'd16611: dataIn1 = 32'd35
; 
32'd16612: dataIn1 = 32'd37
; 
32'd16613: dataIn1 = 32'd48
; 
32'd16614: dataIn1 = 32'd50
; 
32'd16615: dataIn1 = 32'd54
; 
32'd16616: dataIn1 = 32'd58
; 
32'd16617: dataIn1 = 32'd1
; 
32'd16618: dataIn1 = 32'd5
; 
32'd16619: dataIn1 = 32'd9
; 
32'd16620: dataIn1 = 32'd12
; 
32'd16621: dataIn1 = 32'd15
; 
32'd16622: dataIn1 = 32'd16
; 
32'd16623: dataIn1 = 32'd19
; 
32'd16624: dataIn1 = 32'd25
; 
32'd16625: dataIn1 = 32'd31
; 
32'd16626: dataIn1 = 32'd32
; 
32'd16627: dataIn1 = 32'd34
; 
32'd16628: dataIn1 = 32'd36
; 
32'd16629: dataIn1 = 32'd37
; 
32'd16630: dataIn1 = 32'd38
; 
32'd16631: dataIn1 = 32'd41
; 
32'd16632: dataIn1 = 32'd44
; 
32'd16633: dataIn1 = 32'd46
; 
32'd16634: dataIn1 = 32'd49
; 
32'd16635: dataIn1 = 32'd50
; 
32'd16636: dataIn1 = 32'd53
; 
32'd16637: dataIn1 = 32'd56
; 
32'd16638: dataIn1 = 32'd59
; 
32'd16639: dataIn1 = 32'd63
; 
32'd16640: dataIn1 = 32'd5
; 
32'd16641: dataIn1 = 32'd8
; 
32'd16642: dataIn1 = 32'd9
; 
32'd16643: dataIn1 = 32'd10
; 
32'd16644: dataIn1 = 32'd13
; 
32'd16645: dataIn1 = 32'd14
; 
32'd16646: dataIn1 = 32'd22
; 
32'd16647: dataIn1 = 32'd26
; 
32'd16648: dataIn1 = 32'd28
; 
32'd16649: dataIn1 = 32'd29
; 
32'd16650: dataIn1 = 32'd40
; 
32'd16651: dataIn1 = 32'd44
; 
32'd16652: dataIn1 = 32'd45
; 
32'd16653: dataIn1 = 32'd47
; 
32'd16654: dataIn1 = 32'd50
; 
32'd16655: dataIn1 = 32'd58
; 
32'd16656: dataIn1 = 32'd60
; 
32'd16657: dataIn1 = 32'd5
; 
32'd16658: dataIn1 = 32'd6
; 
32'd16659: dataIn1 = 32'd9
; 
32'd16660: dataIn1 = 32'd12
; 
32'd16661: dataIn1 = 32'd14
; 
32'd16662: dataIn1 = 32'd15
; 
32'd16663: dataIn1 = 32'd16
; 
32'd16664: dataIn1 = 32'd19
; 
32'd16665: dataIn1 = 32'd27
; 
32'd16666: dataIn1 = 32'd28
; 
32'd16667: dataIn1 = 32'd31
; 
32'd16668: dataIn1 = 32'd32
; 
32'd16669: dataIn1 = 32'd36
; 
32'd16670: dataIn1 = 32'd41
; 
32'd16671: dataIn1 = 32'd42
; 
32'd16672: dataIn1 = 32'd43
; 
32'd16673: dataIn1 = 32'd46
; 
32'd16674: dataIn1 = 32'd47
; 
32'd16675: dataIn1 = 32'd48
; 
32'd16676: dataIn1 = 32'd49
; 
32'd16677: dataIn1 = 32'd50
; 
32'd16678: dataIn1 = 32'd54
; 
32'd16679: dataIn1 = 32'd56
; 
32'd16680: dataIn1 = 32'd57
; 
32'd16681: dataIn1 = 32'd58
; 
32'd16682: dataIn1 = 32'd62
; 
32'd16683: dataIn1 = 32'd63
; 
32'd16684: dataIn1 = 32'd1
; 
32'd16685: dataIn1 = 32'd3
; 
32'd16686: dataIn1 = 32'd12
; 
32'd16687: dataIn1 = 32'd13
; 
32'd16688: dataIn1 = 32'd14
; 
32'd16689: dataIn1 = 32'd16
; 
32'd16690: dataIn1 = 32'd18
; 
32'd16691: dataIn1 = 32'd23
; 
32'd16692: dataIn1 = 32'd26
; 
32'd16693: dataIn1 = 32'd33
; 
32'd16694: dataIn1 = 32'd34
; 
32'd16695: dataIn1 = 32'd37
; 
32'd16696: dataIn1 = 32'd41
; 
32'd16697: dataIn1 = 32'd44
; 
32'd16698: dataIn1 = 32'd49
; 
32'd16699: dataIn1 = 32'd51
; 
32'd16700: dataIn1 = 32'd52
; 
32'd16701: dataIn1 = 32'd60
; 
32'd16702: dataIn1 = 32'd62
; 
32'd16703: dataIn1 = 32'd5
; 
32'd16704: dataIn1 = 32'd6
; 
32'd16705: dataIn1 = 32'd8
; 
32'd16706: dataIn1 = 32'd12
; 
32'd16707: dataIn1 = 32'd28
; 
32'd16708: dataIn1 = 32'd32
; 
32'd16709: dataIn1 = 32'd33
; 
32'd16710: dataIn1 = 32'd34
; 
32'd16711: dataIn1 = 32'd36
; 
32'd16712: dataIn1 = 32'd37
; 
32'd16713: dataIn1 = 32'd38
; 
32'd16714: dataIn1 = 32'd41
; 
32'd16715: dataIn1 = 32'd46
; 
32'd16716: dataIn1 = 32'd49
; 
32'd16717: dataIn1 = 32'd50
; 
32'd16718: dataIn1 = 32'd52
; 
32'd16719: dataIn1 = 32'd55
; 
32'd16720: dataIn1 = 32'd56
; 
32'd16721: dataIn1 = 32'd57
; 
32'd16722: dataIn1 = 32'd60
; 
32'd16723: dataIn1 = 32'd0
; 
32'd16724: dataIn1 = 32'd1
; 
32'd16725: dataIn1 = 32'd2
; 
32'd16726: dataIn1 = 32'd12
; 
32'd16727: dataIn1 = 32'd17
; 
32'd16728: dataIn1 = 32'd21
; 
32'd16729: dataIn1 = 32'd23
; 
32'd16730: dataIn1 = 32'd25
; 
32'd16731: dataIn1 = 32'd26
; 
32'd16732: dataIn1 = 32'd27
; 
32'd16733: dataIn1 = 32'd29
; 
32'd16734: dataIn1 = 32'd32
; 
32'd16735: dataIn1 = 32'd35
; 
32'd16736: dataIn1 = 32'd37
; 
32'd16737: dataIn1 = 32'd41
; 
32'd16738: dataIn1 = 32'd42
; 
32'd16739: dataIn1 = 32'd46
; 
32'd16740: dataIn1 = 32'd50
; 
32'd16741: dataIn1 = 32'd54
; 
32'd16742: dataIn1 = 32'd55
; 
32'd16743: dataIn1 = 32'd3
; 
32'd16744: dataIn1 = 32'd5
; 
32'd16745: dataIn1 = 32'd7
; 
32'd16746: dataIn1 = 32'd8
; 
32'd16747: dataIn1 = 32'd10
; 
32'd16748: dataIn1 = 32'd11
; 
32'd16749: dataIn1 = 32'd14
; 
32'd16750: dataIn1 = 32'd16
; 
32'd16751: dataIn1 = 32'd17
; 
32'd16752: dataIn1 = 32'd18
; 
32'd16753: dataIn1 = 32'd26
; 
32'd16754: dataIn1 = 32'd27
; 
32'd16755: dataIn1 = 32'd28
; 
32'd16756: dataIn1 = 32'd32
; 
32'd16757: dataIn1 = 32'd33
; 
32'd16758: dataIn1 = 32'd37
; 
32'd16759: dataIn1 = 32'd38
; 
32'd16760: dataIn1 = 32'd50
; 
32'd16761: dataIn1 = 32'd51
; 
32'd16762: dataIn1 = 32'd53
; 
32'd16763: dataIn1 = 32'd60
; 
32'd16764: dataIn1 = 32'd61
; 
32'd16765: dataIn1 = 32'd0
; 
32'd16766: dataIn1 = 32'd5
; 
32'd16767: dataIn1 = 32'd6
; 
32'd16768: dataIn1 = 32'd8
; 
32'd16769: dataIn1 = 32'd11
; 
32'd16770: dataIn1 = 32'd13
; 
32'd16771: dataIn1 = 32'd15
; 
32'd16772: dataIn1 = 32'd17
; 
32'd16773: dataIn1 = 32'd18
; 
32'd16774: dataIn1 = 32'd22
; 
32'd16775: dataIn1 = 32'd23
; 
32'd16776: dataIn1 = 32'd25
; 
32'd16777: dataIn1 = 32'd28
; 
32'd16778: dataIn1 = 32'd35
; 
32'd16779: dataIn1 = 32'd36
; 
32'd16780: dataIn1 = 32'd44
; 
32'd16781: dataIn1 = 32'd45
; 
32'd16782: dataIn1 = 32'd53
; 
32'd16783: dataIn1 = 32'd59
; 
32'd16784: dataIn1 = 32'd60
; 
32'd16785: dataIn1 = 32'd61
; 
32'd16786: dataIn1 = 32'd0
; 
32'd16787: dataIn1 = 32'd2
; 
32'd16788: dataIn1 = 32'd3
; 
32'd16789: dataIn1 = 32'd12
; 
32'd16790: dataIn1 = 32'd17
; 
32'd16791: dataIn1 = 32'd23
; 
32'd16792: dataIn1 = 32'd27
; 
32'd16793: dataIn1 = 32'd30
; 
32'd16794: dataIn1 = 32'd40
; 
32'd16795: dataIn1 = 32'd41
; 
32'd16796: dataIn1 = 32'd43
; 
32'd16797: dataIn1 = 32'd47
; 
32'd16798: dataIn1 = 32'd48
; 
32'd16799: dataIn1 = 32'd53
; 
32'd16800: dataIn1 = 32'd54
; 
32'd16801: dataIn1 = 32'd59
; 
32'd16802: dataIn1 = 32'd0
; 
32'd16803: dataIn1 = 32'd1
; 
32'd16804: dataIn1 = 32'd2
; 
32'd16805: dataIn1 = 32'd3
; 
32'd16806: dataIn1 = 32'd11
; 
32'd16807: dataIn1 = 32'd13
; 
32'd16808: dataIn1 = 32'd14
; 
32'd16809: dataIn1 = 32'd15
; 
32'd16810: dataIn1 = 32'd17
; 
32'd16811: dataIn1 = 32'd19
; 
32'd16812: dataIn1 = 32'd28
; 
32'd16813: dataIn1 = 32'd29
; 
32'd16814: dataIn1 = 32'd31
; 
32'd16815: dataIn1 = 32'd34
; 
32'd16816: dataIn1 = 32'd41
; 
32'd16817: dataIn1 = 32'd47
; 
32'd16818: dataIn1 = 32'd48
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd43; 
32'd3: dataIn2 = 32'd97; 
32'd4: dataIn2 = 32'd13; 
32'd5: dataIn2 = 32'd94; 
32'd6: dataIn2 = 32'd9; 
32'd7: dataIn2 = 32'd83; 
32'd8: dataIn2 = 32'd83; 
32'd9: dataIn2 = 32'd54; 
32'd10: dataIn2 = 32'd92; 
32'd11: dataIn2 = 32'd59; 
32'd12: dataIn2 = 32'd53; 
32'd13: dataIn2 = 32'd83; 
32'd14: dataIn2 = 32'd43; 
32'd15: dataIn2 = 32'd82; 
32'd16: dataIn2 = 32'd67; 
32'd17: dataIn2 = 32'd60; 
32'd18: dataIn2 = 32'd39; 
32'd19: dataIn2 = 32'd9; 
32'd20: dataIn2 = 32'd12; 
32'd21: dataIn2 = 32'd94; 
32'd22: dataIn2 = 32'd89; 
32'd23: dataIn2 = 32'd1; 
32'd24: dataIn2 = 32'd41; 
32'd25: dataIn2 = 32'd49; 
32'd26: dataIn2 = 32'd62; 
32'd27: dataIn2 = 32'd29; 
32'd28: dataIn2 = 32'd0; 
32'd29: dataIn2 = 32'd1; 
32'd30: dataIn2 = 32'd50; 
32'd31: dataIn2 = 32'd80; 
32'd32: dataIn2 = 32'd8; 
32'd33: dataIn2 = 32'd20; 
32'd34: dataIn2 = 32'd10; 
32'd35: dataIn2 = 32'd66; 
32'd36: dataIn2 = 32'd80; 
32'd37: dataIn2 = 32'd56; 
32'd38: dataIn2 = 32'd85; 
32'd39: dataIn2 = 32'd98; 
32'd40: dataIn2 = 32'd8; 
32'd41: dataIn2 = 32'd44; 
32'd42: dataIn2 = 32'd39; 
32'd43: dataIn2 = 32'd76; 
32'd44: dataIn2 = 32'd87; 
32'd45: dataIn2 = 32'd5; 
32'd46: dataIn2 = 32'd45; 
32'd47: dataIn2 = 32'd4; 
32'd48: dataIn2 = 32'd18; 
32'd49: dataIn2 = 32'd2; 
32'd50: dataIn2 = 32'd0; 
32'd51: dataIn2 = 32'd84; 
32'd52: dataIn2 = 32'd50; 
32'd53: dataIn2 = 32'd14; 
32'd54: dataIn2 = 32'd23; 
32'd55: dataIn2 = 32'd26; 
32'd56: dataIn2 = 32'd6; 
32'd57: dataIn2 = 32'd68; 
32'd58: dataIn2 = 32'd30; 
32'd59: dataIn2 = 32'd47; 
32'd60: dataIn2 = 32'd42; 
32'd61: dataIn2 = 32'd52; 
32'd62: dataIn2 = 32'd29; 
32'd63: dataIn2 = 32'd5; 
32'd64: dataIn2 = 32'd57; 
32'd65: dataIn2 = 32'd39; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd330: dataIn2 = 32'd18; 
32'd331: dataIn2 = 32'd5; 
32'd332: dataIn2 = 32'd49; 
32'd333: dataIn2 = 32'd72; 
32'd334: dataIn2 = 32'd19; 
32'd335: dataIn2 = 32'd34; 
32'd336: dataIn2 = 32'd53; 
32'd337: dataIn2 = 32'd49; 
32'd338: dataIn2 = 32'd79; 
32'd339: dataIn2 = 32'd7; 
32'd340: dataIn2 = 32'd35; 
32'd341: dataIn2 = 32'd87; 
32'd342: dataIn2 = 32'd0; 
32'd343: dataIn2 = 32'd89; 
32'd344: dataIn2 = 32'd95; 
32'd345: dataIn2 = 32'd66; 
32'd346: dataIn2 = 32'd83; 
32'd347: dataIn2 = 32'd95; 
32'd348: dataIn2 = 32'd11; 
32'd349: dataIn2 = 32'd9; 
32'd350: dataIn2 = 32'd37; 
32'd351: dataIn2 = 32'd21; 
32'd352: dataIn2 = 32'd41; 
32'd353: dataIn2 = 32'd86; 
32'd354: dataIn2 = 32'd99; 
32'd355: dataIn2 = 32'd91; 
32'd356: dataIn2 = 32'd10; 
32'd357: dataIn2 = 32'd93; 
32'd358: dataIn2 = 32'd71; 
32'd359: dataIn2 = 32'd44; 
32'd360: dataIn2 = 32'd81; 
32'd361: dataIn2 = 32'd26; 
32'd362: dataIn2 = 32'd65; 
32'd363: dataIn2 = 32'd97; 
32'd364: dataIn2 = 32'd31; 
32'd365: dataIn2 = 32'd64; 
32'd366: dataIn2 = 32'd67; 
32'd367: dataIn2 = 32'd85; 
32'd368: dataIn2 = 32'd45; 
32'd369: dataIn2 = 32'd78; 
32'd370: dataIn2 = 32'd100; 
32'd371: dataIn2 = 32'd89; 
32'd372: dataIn2 = 32'd32; 
32'd373: dataIn2 = 32'd8; 
32'd374: dataIn2 = 32'd93; 
32'd375: dataIn2 = 32'd65; 
32'd376: dataIn2 = 32'd26; 
32'd377: dataIn2 = 32'd100; 
32'd378: dataIn2 = 32'd89; 
32'd379: dataIn2 = 32'd62; 
32'd380: dataIn2 = 32'd81; 
32'd381: dataIn2 = 32'd97; 
32'd382: dataIn2 = 32'd37; 
32'd383: dataIn2 = 32'd54; 
32'd384: dataIn2 = 32'd87; 
32'd385: dataIn2 = 32'd51; 
32'd386: dataIn2 = 32'd74; 
32'd387: dataIn2 = 32'd45; 
32'd388: dataIn2 = 32'd61; 
32'd389: dataIn2 = 32'd20; 
32'd390: dataIn2 = 32'd87; 
32'd391: dataIn2 = 32'd91; 
32'd392: dataIn2 = 32'd39; 
32'd393: dataIn2 = 32'd68; 
32'd394: dataIn2 = 32'd65; 
32'd395: dataIn2 = 32'd19; 
32'd396: dataIn2 = 32'd66; 
32'd397: dataIn2 = 32'd49; 
32'd398: dataIn2 = 32'd94; 
32'd399: dataIn2 = 32'd71; 
32'd400: dataIn2 = 32'd94; 
32'd401: dataIn2 = 32'd29; 
32'd402: dataIn2 = 32'd67; 
32'd403: dataIn2 = 32'd67; 
32'd404: dataIn2 = 32'd43; 
32'd405: dataIn2 = 32'd22; 
32'd406: dataIn2 = 32'd14; 
32'd407: dataIn2 = 32'd64; 
32'd408: dataIn2 = 32'd19; 
32'd409: dataIn2 = 32'd11; 
32'd410: dataIn2 = 32'd69; 
32'd411: dataIn2 = 32'd92; 
32'd412: dataIn2 = 32'd65; 
32'd413: dataIn2 = 32'd92; 
32'd414: dataIn2 = 32'd48; 
32'd415: dataIn2 = 32'd25; 
32'd416: dataIn2 = 32'd44; 
32'd417: dataIn2 = 32'd22; 
32'd418: dataIn2 = 32'd13; 
32'd419: dataIn2 = 32'd62; 
32'd420: dataIn2 = 32'd32; 
32'd421: dataIn2 = 32'd5; 
32'd422: dataIn2 = 32'd42; 
32'd423: dataIn2 = 32'd77; 
32'd424: dataIn2 = 32'd91; 
32'd425: dataIn2 = 32'd98; 
32'd426: dataIn2 = 32'd13; 
32'd427: dataIn2 = 32'd12; 
32'd428: dataIn2 = 32'd44; 
32'd429: dataIn2 = 32'd93; 
32'd430: dataIn2 = 32'd100; 
32'd431: dataIn2 = 32'd57; 
32'd432: dataIn2 = 32'd61; 
32'd433: dataIn2 = 32'd58; 
32'd434: dataIn2 = 32'd56; 
32'd435: dataIn2 = 32'd66; 
32'd436: dataIn2 = 32'd17; 
32'd437: dataIn2 = 32'd62; 
32'd438: dataIn2 = 32'd54; 
32'd439: dataIn2 = 32'd16; 
32'd440: dataIn2 = 32'd39; 
32'd441: dataIn2 = 32'd67; 
32'd442: dataIn2 = 32'd13; 
32'd443: dataIn2 = 32'd65; 
32'd444: dataIn2 = 32'd77; 
32'd445: dataIn2 = 32'd22; 
32'd446: dataIn2 = 32'd12; 
32'd447: dataIn2 = 32'd46; 
32'd448: dataIn2 = 32'd13; 
32'd449: dataIn2 = 32'd10; 
32'd450: dataIn2 = 32'd96; 
32'd451: dataIn2 = 32'd80; 
32'd452: dataIn2 = 32'd61; 
32'd453: dataIn2 = 32'd49; 
32'd454: dataIn2 = 32'd81; 
32'd455: dataIn2 = 32'd49; 
32'd456: dataIn2 = 32'd98; 
32'd457: dataIn2 = 32'd63; 
32'd458: dataIn2 = 32'd59; 
32'd459: dataIn2 = 32'd32; 
32'd460: dataIn2 = 32'd76; 
32'd461: dataIn2 = 32'd70; 
32'd462: dataIn2 = 32'd14; 
32'd463: dataIn2 = 32'd39; 
32'd464: dataIn2 = 32'd14; 
32'd465: dataIn2 = 32'd13; 
32'd466: dataIn2 = 32'd84; 
32'd467: dataIn2 = 32'd11; 
32'd468: dataIn2 = 32'd62; 
32'd469: dataIn2 = 32'd67; 
32'd470: dataIn2 = 32'd3; 
32'd471: dataIn2 = 32'd38; 
32'd472: dataIn2 = 32'd87; 
32'd473: dataIn2 = 32'd65; 
32'd474: dataIn2 = 32'd93; 
32'd475: dataIn2 = 32'd35; 
32'd476: dataIn2 = 32'd12; 
32'd477: dataIn2 = 32'd53; 
32'd478: dataIn2 = 32'd27; 
32'd479: dataIn2 = 32'd51; 
32'd480: dataIn2 = 32'd27; 
32'd481: dataIn2 = 32'd31; 
32'd482: dataIn2 = 32'd97; 
32'd483: dataIn2 = 32'd4; 
32'd484: dataIn2 = 32'd37; 
32'd485: dataIn2 = 32'd22; 
32'd486: dataIn2 = 32'd68; 
32'd487: dataIn2 = 32'd41; 
32'd488: dataIn2 = 32'd36; 
32'd489: dataIn2 = 32'd53; 
32'd490: dataIn2 = 32'd65; 
32'd491: dataIn2 = 32'd64; 
32'd492: dataIn2 = 32'd81; 
32'd493: dataIn2 = 32'd91; 
32'd494: dataIn2 = 32'd100; 
32'd495: dataIn2 = 32'd14; 
32'd496: dataIn2 = 32'd19; 
32'd497: dataIn2 = 32'd21; 
32'd498: dataIn2 = 32'd13; 
32'd499: dataIn2 = 32'd6; 
32'd500: dataIn2 = 32'd25; 
32'd501: dataIn2 = 32'd26; 
32'd502: dataIn2 = 32'd25; 
32'd503: dataIn2 = 32'd64; 
32'd504: dataIn2 = 32'd3; 
32'd505: dataIn2 = 32'd45; 
32'd506: dataIn2 = 32'd76; 
32'd507: dataIn2 = 32'd90; 
32'd508: dataIn2 = 32'd95; 
32'd509: dataIn2 = 32'd45; 
32'd510: dataIn2 = 32'd23; 
32'd511: dataIn2 = 32'd40; 
32'd512: dataIn2 = 32'd31; 
32'd513: dataIn2 = 32'd18; 
32'd514: dataIn2 = 32'd8; 
32'd515: dataIn2 = 32'd5; 
32'd516: dataIn2 = 32'd88; 
32'd517: dataIn2 = 32'd51; 
32'd518: dataIn2 = 32'd6; 
32'd519: dataIn2 = 32'd33; 
32'd520: dataIn2 = 32'd13; 
32'd521: dataIn2 = 32'd32; 
32'd522: dataIn2 = 32'd63; 
32'd523: dataIn2 = 32'd9; 
32'd524: dataIn2 = 32'd77; 
32'd525: dataIn2 = 32'd98; 
32'd526: dataIn2 = 32'd17; 
32'd527: dataIn2 = 32'd8; 
32'd528: dataIn2 = 32'd84; 
32'd529: dataIn2 = 32'd90; 
32'd530: dataIn2 = 32'd6; 
32'd531: dataIn2 = 32'd45; 
32'd532: dataIn2 = 32'd31; 
32'd533: dataIn2 = 32'd43; 
32'd534: dataIn2 = 32'd9; 
32'd535: dataIn2 = 32'd23; 
32'd536: dataIn2 = 32'd9; 
32'd537: dataIn2 = 32'd37; 
32'd538: dataIn2 = 32'd12; 
32'd539: dataIn2 = 32'd96; 
32'd540: dataIn2 = 32'd83; 
32'd541: dataIn2 = 32'd72; 
32'd542: dataIn2 = 32'd98; 
32'd543: dataIn2 = 32'd39; 
32'd544: dataIn2 = 32'd29; 
32'd545: dataIn2 = 32'd75; 
32'd546: dataIn2 = 32'd16; 
32'd547: dataIn2 = 32'd87; 
32'd548: dataIn2 = 32'd68; 
32'd549: dataIn2 = 32'd87; 
32'd550: dataIn2 = 32'd29; 
32'd551: dataIn2 = 32'd98; 
32'd552: dataIn2 = 32'd3; 
32'd553: dataIn2 = 32'd37; 
32'd554: dataIn2 = 32'd41; 
32'd555: dataIn2 = 32'd12; 
32'd556: dataIn2 = 32'd74; 
32'd557: dataIn2 = 32'd87; 
32'd558: dataIn2 = 32'd45; 
32'd559: dataIn2 = 32'd35; 
32'd560: dataIn2 = 32'd74; 
32'd561: dataIn2 = 32'd3; 
32'd562: dataIn2 = 32'd74; 
32'd563: dataIn2 = 32'd99; 
32'd564: dataIn2 = 32'd81; 
32'd565: dataIn2 = 32'd75; 
32'd566: dataIn2 = 32'd65; 
32'd567: dataIn2 = 32'd79; 
32'd568: dataIn2 = 32'd78; 
32'd569: dataIn2 = 32'd52; 
32'd570: dataIn2 = 32'd30; 
32'd571: dataIn2 = 32'd52; 
32'd572: dataIn2 = 32'd67; 
32'd573: dataIn2 = 32'd13; 
32'd574: dataIn2 = 32'd34; 
32'd575: dataIn2 = 32'd14; 
32'd576: dataIn2 = 32'd22; 
32'd577: dataIn2 = 32'd32; 
32'd578: dataIn2 = 32'd13; 
32'd579: dataIn2 = 32'd17; 
32'd580: dataIn2 = 32'd95; 
32'd581: dataIn2 = 32'd4; 
32'd582: dataIn2 = 32'd8; 
32'd583: dataIn2 = 32'd62; 
32'd584: dataIn2 = 32'd54; 
32'd585: dataIn2 = 32'd32; 
32'd586: dataIn2 = 32'd54; 
32'd587: dataIn2 = 32'd82; 
32'd588: dataIn2 = 32'd85; 
32'd589: dataIn2 = 32'd39; 
32'd590: dataIn2 = 32'd74; 
32'd591: dataIn2 = 32'd89; 
32'd592: dataIn2 = 32'd65; 
32'd593: dataIn2 = 32'd48; 
32'd594: dataIn2 = 32'd88; 
32'd595: dataIn2 = 32'd90; 
32'd596: dataIn2 = 32'd12; 
32'd597: dataIn2 = 32'd63; 
32'd598: dataIn2 = 32'd17; 
32'd599: dataIn2 = 32'd35; 
32'd600: dataIn2 = 32'd78; 
32'd601: dataIn2 = 32'd68; 
32'd602: dataIn2 = 32'd58; 
32'd603: dataIn2 = 32'd17; 
32'd604: dataIn2 = 32'd27; 
32'd605: dataIn2 = 32'd36; 
32'd606: dataIn2 = 32'd3; 
32'd607: dataIn2 = 32'd5; 
32'd608: dataIn2 = 32'd19; 
32'd609: dataIn2 = 32'd83; 
32'd610: dataIn2 = 32'd93; 
32'd611: dataIn2 = 32'd37; 
32'd612: dataIn2 = 32'd31; 
32'd613: dataIn2 = 32'd54; 
32'd614: dataIn2 = 32'd29; 
32'd615: dataIn2 = 32'd24; 
32'd616: dataIn2 = 32'd96; 
32'd617: dataIn2 = 32'd7; 
32'd618: dataIn2 = 32'd69; 
32'd619: dataIn2 = 32'd69; 
32'd620: dataIn2 = 32'd14; 
32'd621: dataIn2 = 32'd55; 
32'd622: dataIn2 = 32'd11; 
32'd623: dataIn2 = 32'd13; 
32'd624: dataIn2 = 32'd87; 
32'd625: dataIn2 = 32'd64; 
32'd626: dataIn2 = 32'd71; 
32'd627: dataIn2 = 32'd40; 
32'd628: dataIn2 = 32'd21; 
32'd629: dataIn2 = 32'd2; 
32'd630: dataIn2 = 32'd69; 
32'd631: dataIn2 = 32'd42; 
32'd632: dataIn2 = 32'd16; 
32'd633: dataIn2 = 32'd45; 
32'd634: dataIn2 = 32'd0; 
32'd635: dataIn2 = 32'd71; 
32'd636: dataIn2 = 32'd78; 
32'd637: dataIn2 = 32'd12; 
32'd638: dataIn2 = 32'd15; 
32'd639: dataIn2 = 32'd87; 
32'd640: dataIn2 = 32'd93; 
32'd641: dataIn2 = 32'd21; 
32'd642: dataIn2 = 32'd72; 
32'd643: dataIn2 = 32'd20; 
32'd644: dataIn2 = 32'd73; 
32'd645: dataIn2 = 32'd90; 
32'd646: dataIn2 = 32'd40; 
32'd647: dataIn2 = 32'd10; 
32'd648: dataIn2 = 32'd73; 
32'd649: dataIn2 = 32'd60; 
32'd650: dataIn2 = 32'd3; 
32'd651: dataIn2 = 32'd15; 
32'd652: dataIn2 = 32'd53; 
32'd653: dataIn2 = 32'd89; 
32'd654: dataIn2 = 32'd11; 
32'd655: dataIn2 = 32'd93; 
32'd656: dataIn2 = 32'd54; 
32'd657: dataIn2 = 32'd88; 
32'd658: dataIn2 = 32'd33; 
32'd659: dataIn2 = 32'd57; 
32'd660: dataIn2 = 32'd92; 
32'd661: dataIn2 = 32'd43; 
32'd662: dataIn2 = 32'd78; 
32'd663: dataIn2 = 32'd80; 
32'd664: dataIn2 = 32'd63; 
32'd665: dataIn2 = 32'd30; 
32'd666: dataIn2 = 32'd90; 
32'd667: dataIn2 = 32'd69; 
32'd668: dataIn2 = 32'd82; 
32'd669: dataIn2 = 32'd94; 
32'd670: dataIn2 = 32'd53; 
32'd671: dataIn2 = 32'd8; 
32'd672: dataIn2 = 32'd23; 
32'd673: dataIn2 = 32'd22; 
32'd674: dataIn2 = 32'd25; 
32'd675: dataIn2 = 32'd83; 
32'd676: dataIn2 = 32'd89; 
32'd677: dataIn2 = 32'd68; 
32'd678: dataIn2 = 32'd75; 
32'd679: dataIn2 = 32'd5; 
32'd680: dataIn2 = 32'd55; 
32'd681: dataIn2 = 32'd18; 
32'd682: dataIn2 = 32'd97; 
32'd683: dataIn2 = 32'd91; 
32'd684: dataIn2 = 32'd24; 
32'd685: dataIn2 = 32'd11; 
32'd686: dataIn2 = 32'd96; 
32'd687: dataIn2 = 32'd79; 
32'd688: dataIn2 = 32'd63; 
32'd689: dataIn2 = 32'd62; 
32'd690: dataIn2 = 32'd6; 
32'd691: dataIn2 = 32'd27; 
32'd692: dataIn2 = 32'd9; 
32'd693: dataIn2 = 32'd59; 
32'd694: dataIn2 = 32'd41; 
32'd695: dataIn2 = 32'd86; 
32'd696: dataIn2 = 32'd29; 
32'd697: dataIn2 = 32'd75; 
32'd698: dataIn2 = 32'd10; 
32'd699: dataIn2 = 32'd18; 
32'd700: dataIn2 = 32'd88; 
32'd701: dataIn2 = 32'd41; 
32'd702: dataIn2 = 32'd66; 
32'd703: dataIn2 = 32'd60; 
32'd704: dataIn2 = 32'd32; 
32'd705: dataIn2 = 32'd22; 
32'd706: dataIn2 = 32'd31; 
32'd707: dataIn2 = 32'd36; 
32'd708: dataIn2 = 32'd77; 
32'd709: dataIn2 = 32'd67; 
32'd710: dataIn2 = 32'd76; 
32'd711: dataIn2 = 32'd51; 
32'd712: dataIn2 = 32'd54; 
32'd713: dataIn2 = 32'd20; 
32'd714: dataIn2 = 32'd14; 
32'd715: dataIn2 = 32'd59; 
32'd716: dataIn2 = 32'd7; 
32'd717: dataIn2 = 32'd11; 
32'd718: dataIn2 = 32'd32; 
32'd719: dataIn2 = 32'd43; 
32'd720: dataIn2 = 32'd85; 
32'd721: dataIn2 = 32'd48; 
32'd722: dataIn2 = 32'd15; 
32'd723: dataIn2 = 32'd10; 
32'd724: dataIn2 = 32'd76; 
32'd725: dataIn2 = 32'd68; 
32'd726: dataIn2 = 32'd47; 
32'd727: dataIn2 = 32'd67; 
32'd728: dataIn2 = 32'd20; 
32'd729: dataIn2 = 32'd75; 
32'd730: dataIn2 = 32'd52; 
32'd731: dataIn2 = 32'd84; 
32'd732: dataIn2 = 32'd85; 
32'd733: dataIn2 = 32'd3; 
32'd734: dataIn2 = 32'd50; 
32'd735: dataIn2 = 32'd45; 
32'd736: dataIn2 = 32'd46; 
32'd737: dataIn2 = 32'd22; 
32'd738: dataIn2 = 32'd11; 
32'd739: dataIn2 = 32'd21; 
32'd740: dataIn2 = 32'd95; 
32'd741: dataIn2 = 32'd97; 
32'd742: dataIn2 = 32'd15; 
32'd743: dataIn2 = 32'd57; 
32'd744: dataIn2 = 32'd31; 
32'd745: dataIn2 = 32'd39; 
32'd746: dataIn2 = 32'd89; 
32'd747: dataIn2 = 32'd97; 
32'd748: dataIn2 = 32'd46; 
32'd749: dataIn2 = 32'd79; 
32'd750: dataIn2 = 32'd75; 
32'd751: dataIn2 = 32'd2; 
32'd752: dataIn2 = 32'd16; 
32'd753: dataIn2 = 32'd96; 
32'd754: dataIn2 = 32'd59; 
32'd755: dataIn2 = 32'd24; 
32'd756: dataIn2 = 32'd29; 
32'd757: dataIn2 = 32'd98; 
32'd758: dataIn2 = 32'd71; 
32'd759: dataIn2 = 32'd35; 
32'd760: dataIn2 = 32'd13; 
32'd761: dataIn2 = 32'd29; 
32'd762: dataIn2 = 32'd23; 
32'd763: dataIn2 = 32'd64; 
32'd764: dataIn2 = 32'd15; 
32'd765: dataIn2 = 32'd87; 
32'd766: dataIn2 = 32'd48; 
32'd767: dataIn2 = 32'd29; 
32'd768: dataIn2 = 32'd55; 
32'd769: dataIn2 = 32'd59; 
32'd770: dataIn2 = 32'd92; 
32'd771: dataIn2 = 32'd30; 
32'd772: dataIn2 = 32'd54; 
32'd773: dataIn2 = 32'd36; 
32'd774: dataIn2 = 32'd24; 
32'd775: dataIn2 = 32'd76; 
32'd776: dataIn2 = 32'd48; 
32'd777: dataIn2 = 32'd18; 
32'd778: dataIn2 = 32'd35; 
32'd779: dataIn2 = 32'd75; 
32'd780: dataIn2 = 32'd45; 
32'd781: dataIn2 = 32'd86; 
32'd782: dataIn2 = 32'd84; 
32'd783: dataIn2 = 32'd45; 
32'd784: dataIn2 = 32'd100; 
32'd785: dataIn2 = 32'd65; 
32'd786: dataIn2 = 32'd76; 
32'd787: dataIn2 = 32'd80; 
32'd788: dataIn2 = 32'd39; 
32'd789: dataIn2 = 32'd1; 
32'd790: dataIn2 = 32'd47; 
32'd791: dataIn2 = 32'd1; 
32'd792: dataIn2 = 32'd61; 
32'd793: dataIn2 = 32'd63; 
32'd794: dataIn2 = 32'd58; 
32'd795: dataIn2 = 32'd46; 
32'd796: dataIn2 = 32'd72; 
32'd797: dataIn2 = 32'd95; 
32'd798: dataIn2 = 32'd37; 
32'd799: dataIn2 = 32'd13; 
32'd800: dataIn2 = 32'd17; 
32'd801: dataIn2 = 32'd35; 
32'd802: dataIn2 = 32'd29; 
32'd803: dataIn2 = 32'd63; 
32'd804: dataIn2 = 32'd22; 
32'd805: dataIn2 = 32'd45; 
32'd806: dataIn2 = 32'd54; 
32'd807: dataIn2 = 32'd33; 
32'd808: dataIn2 = 32'd27; 
32'd809: dataIn2 = 32'd42; 
32'd810: dataIn2 = 32'd34; 
32'd811: dataIn2 = 32'd96; 
32'd812: dataIn2 = 32'd13; 
32'd813: dataIn2 = 32'd6; 
32'd814: dataIn2 = 32'd83; 
32'd815: dataIn2 = 32'd50; 
32'd816: dataIn2 = 32'd15; 
32'd817: dataIn2 = 32'd30; 
32'd818: dataIn2 = 32'd41; 
32'd819: dataIn2 = 32'd15; 
32'd820: dataIn2 = 32'd54; 
32'd821: dataIn2 = 32'd69; 
32'd822: dataIn2 = 32'd70; 
32'd823: dataIn2 = 32'd83; 
32'd824: dataIn2 = 32'd19; 
32'd825: dataIn2 = 32'd21; 
32'd826: dataIn2 = 32'd3; 
32'd827: dataIn2 = 32'd69; 
32'd828: dataIn2 = 32'd91; 
32'd829: dataIn2 = 32'd43; 
32'd830: dataIn2 = 32'd18; 
32'd831: dataIn2 = 32'd91; 
32'd832: dataIn2 = 32'd55; 
32'd833: dataIn2 = 32'd16; 
32'd834: dataIn2 = 32'd44; 
32'd835: dataIn2 = 32'd79; 
32'd836: dataIn2 = 32'd12; 
32'd837: dataIn2 = 32'd28; 
32'd838: dataIn2 = 32'd8; 
32'd839: dataIn2 = 32'd99; 
32'd840: dataIn2 = 32'd26; 
32'd841: dataIn2 = 32'd80; 
32'd842: dataIn2 = 32'd96; 
32'd843: dataIn2 = 32'd23; 
32'd844: dataIn2 = 32'd53; 
32'd845: dataIn2 = 32'd45; 
32'd846: dataIn2 = 32'd51; 
32'd847: dataIn2 = 32'd44; 
32'd848: dataIn2 = 32'd83; 
32'd849: dataIn2 = 32'd69; 
32'd850: dataIn2 = 32'd21; 
32'd851: dataIn2 = 32'd22; 
32'd852: dataIn2 = 32'd66; 
32'd853: dataIn2 = 32'd47; 
32'd854: dataIn2 = 32'd39; 
32'd855: dataIn2 = 32'd0; 
32'd856: dataIn2 = 32'd49; 
32'd857: dataIn2 = 32'd23; 
32'd858: dataIn2 = 32'd47; 
32'd859: dataIn2 = 32'd72; 
32'd860: dataIn2 = 32'd54; 
32'd861: dataIn2 = 32'd39; 
32'd862: dataIn2 = 32'd63; 
32'd863: dataIn2 = 32'd88; 
32'd864: dataIn2 = 32'd67; 
32'd865: dataIn2 = 32'd6; 
32'd866: dataIn2 = 32'd83; 
32'd867: dataIn2 = 32'd59; 
32'd868: dataIn2 = 32'd22; 
32'd869: dataIn2 = 32'd55; 
32'd870: dataIn2 = 32'd4; 
32'd871: dataIn2 = 32'd81; 
32'd872: dataIn2 = 32'd2; 
32'd873: dataIn2 = 32'd38; 
32'd874: dataIn2 = 32'd33; 
32'd875: dataIn2 = 32'd47; 
32'd876: dataIn2 = 32'd45; 
32'd877: dataIn2 = 32'd62; 
32'd878: dataIn2 = 32'd61; 
32'd879: dataIn2 = 32'd13; 
32'd880: dataIn2 = 32'd87; 
32'd881: dataIn2 = 32'd54; 
32'd882: dataIn2 = 32'd41; 
32'd883: dataIn2 = 32'd73; 
32'd884: dataIn2 = 32'd25; 
32'd885: dataIn2 = 32'd68; 
32'd886: dataIn2 = 32'd58; 
32'd887: dataIn2 = 32'd61; 
32'd888: dataIn2 = 32'd53; 
32'd889: dataIn2 = 32'd8; 
32'd890: dataIn2 = 32'd10; 
32'd891: dataIn2 = 32'd81; 
32'd892: dataIn2 = 32'd96; 
32'd893: dataIn2 = 32'd71; 
32'd894: dataIn2 = 32'd38; 
32'd895: dataIn2 = 32'd91; 
32'd896: dataIn2 = 32'd17; 
32'd897: dataIn2 = 32'd8; 
32'd898: dataIn2 = 32'd77; 
32'd899: dataIn2 = 32'd37; 
32'd900: dataIn2 = 32'd46; 
32'd901: dataIn2 = 32'd25; 
32'd902: dataIn2 = 32'd64; 
32'd903: dataIn2 = 32'd7; 
32'd904: dataIn2 = 32'd92; 
32'd905: dataIn2 = 32'd44; 
32'd906: dataIn2 = 32'd61; 
32'd907: dataIn2 = 32'd49; 
32'd908: dataIn2 = 32'd88; 
32'd909: dataIn2 = 32'd30; 
32'd910: dataIn2 = 32'd24; 
32'd911: dataIn2 = 32'd88; 
32'd912: dataIn2 = 32'd63; 
32'd913: dataIn2 = 32'd43; 
32'd914: dataIn2 = 32'd17; 
32'd915: dataIn2 = 32'd7; 
32'd916: dataIn2 = 32'd24; 
32'd917: dataIn2 = 32'd60; 
32'd918: dataIn2 = 32'd71; 
32'd919: dataIn2 = 32'd89; 
32'd920: dataIn2 = 32'd9; 
32'd921: dataIn2 = 32'd6; 
32'd922: dataIn2 = 32'd18; 
32'd923: dataIn2 = 32'd68; 
32'd924: dataIn2 = 32'd56; 
32'd925: dataIn2 = 32'd24; 
32'd926: dataIn2 = 32'd25; 
32'd927: dataIn2 = 32'd12; 
32'd928: dataIn2 = 32'd69; 
32'd929: dataIn2 = 32'd24; 
32'd930: dataIn2 = 32'd37; 
32'd931: dataIn2 = 32'd61; 
32'd932: dataIn2 = 32'd91; 
32'd933: dataIn2 = 32'd38; 
32'd934: dataIn2 = 32'd63; 
32'd935: dataIn2 = 32'd31; 
32'd936: dataIn2 = 32'd91; 
32'd937: dataIn2 = 32'd69; 
32'd938: dataIn2 = 32'd63; 
32'd939: dataIn2 = 32'd62; 
32'd940: dataIn2 = 32'd69; 
32'd941: dataIn2 = 32'd13; 
32'd942: dataIn2 = 32'd67; 
32'd943: dataIn2 = 32'd14; 
32'd944: dataIn2 = 32'd15; 
32'd945: dataIn2 = 32'd84; 
32'd946: dataIn2 = 32'd33; 
32'd947: dataIn2 = 32'd22; 
32'd948: dataIn2 = 32'd91; 
32'd949: dataIn2 = 32'd84; 
32'd950: dataIn2 = 32'd61; 
32'd951: dataIn2 = 32'd54; 
32'd952: dataIn2 = 32'd30; 
32'd953: dataIn2 = 32'd85; 
32'd954: dataIn2 = 32'd83; 
32'd955: dataIn2 = 32'd4; 
32'd956: dataIn2 = 32'd84; 
32'd957: dataIn2 = 32'd2; 
32'd958: dataIn2 = 32'd29; 
32'd959: dataIn2 = 32'd60; 
32'd960: dataIn2 = 32'd67; 
32'd961: dataIn2 = 32'd87; 
32'd962: dataIn2 = 32'd30; 
32'd963: dataIn2 = 32'd65; 
32'd964: dataIn2 = 32'd95; 
32'd965: dataIn2 = 32'd2; 
32'd966: dataIn2 = 32'd5; 
32'd967: dataIn2 = 32'd78; 
32'd968: dataIn2 = 32'd13; 
32'd969: dataIn2 = 32'd14; 
32'd970: dataIn2 = 32'd45; 
32'd971: dataIn2 = 32'd49; 
32'd972: dataIn2 = 32'd86; 
32'd973: dataIn2 = 32'd54; 
32'd974: dataIn2 = 32'd39; 
32'd975: dataIn2 = 32'd68; 
32'd976: dataIn2 = 32'd23; 
32'd977: dataIn2 = 32'd62; 
32'd978: dataIn2 = 32'd89; 
32'd979: dataIn2 = 32'd30; 
32'd980: dataIn2 = 32'd58; 
32'd981: dataIn2 = 32'd31; 
32'd982: dataIn2 = 32'd5; 
32'd983: dataIn2 = 32'd3; 
32'd984: dataIn2 = 32'd55; 
32'd985: dataIn2 = 32'd52; 
32'd986: dataIn2 = 32'd59; 
32'd987: dataIn2 = 32'd88; 
32'd988: dataIn2 = 32'd7; 
32'd989: dataIn2 = 32'd5; 
32'd990: dataIn2 = 32'd53; 
32'd991: dataIn2 = 32'd25; 
32'd992: dataIn2 = 32'd10; 
32'd993: dataIn2 = 32'd10; 
32'd994: dataIn2 = 32'd75; 
32'd995: dataIn2 = 32'd77; 
32'd996: dataIn2 = 32'd80; 
32'd997: dataIn2 = 32'd91; 
32'd998: dataIn2 = 32'd54; 
32'd999: dataIn2 = 32'd97; 
32'd1000: dataIn2 = 32'd61; 
32'd1001: dataIn2 = 32'd21; 
32'd1002: dataIn2 = 32'd43; 
32'd1003: dataIn2 = 32'd31; 
32'd1004: dataIn2 = 32'd89; 
32'd1005: dataIn2 = 32'd52; 
32'd1006: dataIn2 = 32'd75; 
32'd1007: dataIn2 = 32'd27; 
32'd1008: dataIn2 = 32'd90; 
32'd1009: dataIn2 = 32'd74; 
32'd1010: dataIn2 = 32'd33; 
32'd1011: dataIn2 = 32'd80; 
32'd1012: dataIn2 = 32'd18; 
32'd1013: dataIn2 = 32'd99; 
32'd1014: dataIn2 = 32'd89; 
32'd1015: dataIn2 = 32'd73; 
32'd1016: dataIn2 = 32'd52; 
32'd1017: dataIn2 = 32'd88; 
32'd1018: dataIn2 = 32'd72; 
32'd1019: dataIn2 = 32'd92; 
32'd1020: dataIn2 = 32'd92; 
32'd1021: dataIn2 = 32'd43; 
32'd1022: dataIn2 = 32'd44; 
32'd1023: dataIn2 = 32'd80; 
32'd1024: dataIn2 = 32'd39; 
32'd1025: dataIn2 = 32'd49; 
32'd1026: dataIn2 = 32'd5; 
32'd1027: dataIn2 = 32'd93; 
32'd1028: dataIn2 = 32'd41; 
32'd1029: dataIn2 = 32'd27; 
32'd1030: dataIn2 = 32'd14; 
32'd1031: dataIn2 = 32'd60; 
32'd1032: dataIn2 = 32'd43; 
32'd1033: dataIn2 = 32'd67; 
32'd1034: dataIn2 = 32'd17; 
32'd1035: dataIn2 = 32'd89; 
32'd1036: dataIn2 = 32'd3; 
32'd1037: dataIn2 = 32'd98; 
32'd1038: dataIn2 = 32'd23; 
32'd1039: dataIn2 = 32'd91; 
32'd1040: dataIn2 = 32'd51; 
32'd1041: dataIn2 = 32'd53; 
32'd1042: dataIn2 = 32'd35; 
32'd1043: dataIn2 = 32'd73; 
32'd1044: dataIn2 = 32'd52; 
32'd1045: dataIn2 = 32'd38; 
32'd1046: dataIn2 = 32'd60; 
32'd1047: dataIn2 = 32'd18; 
32'd1048: dataIn2 = 32'd11; 
32'd1049: dataIn2 = 32'd78; 
32'd1050: dataIn2 = 32'd81; 
32'd1051: dataIn2 = 32'd89; 
32'd1052: dataIn2 = 32'd13; 
32'd1053: dataIn2 = 32'd14; 
32'd1054: dataIn2 = 32'd15; 
32'd1055: dataIn2 = 32'd0; 
32'd1056: dataIn2 = 32'd94; 
32'd1057: dataIn2 = 32'd2; 
32'd1058: dataIn2 = 32'd61; 
32'd1059: dataIn2 = 32'd61; 
32'd1060: dataIn2 = 32'd70; 
32'd1061: dataIn2 = 32'd50; 
32'd1062: dataIn2 = 32'd67; 
32'd1063: dataIn2 = 32'd29; 
32'd1064: dataIn2 = 32'd8; 
32'd1065: dataIn2 = 32'd36; 
32'd1066: dataIn2 = 32'd66; 
32'd1067: dataIn2 = 32'd50; 
32'd1068: dataIn2 = 32'd39; 
32'd1069: dataIn2 = 32'd100; 
32'd1070: dataIn2 = 32'd56; 
32'd1071: dataIn2 = 32'd9; 
32'd1072: dataIn2 = 32'd34; 
32'd1073: dataIn2 = 32'd98; 
32'd1074: dataIn2 = 32'd46; 
32'd1075: dataIn2 = 32'd18; 
32'd1076: dataIn2 = 32'd80; 
32'd1077: dataIn2 = 32'd24; 
32'd1078: dataIn2 = 32'd15; 
32'd1079: dataIn2 = 32'd3; 
32'd1080: dataIn2 = 32'd74; 
32'd1081: dataIn2 = 32'd90; 
32'd1082: dataIn2 = 32'd0; 
32'd1083: dataIn2 = 32'd79; 
32'd1084: dataIn2 = 32'd15; 
32'd1085: dataIn2 = 32'd51; 
32'd1086: dataIn2 = 32'd78; 
32'd1087: dataIn2 = 32'd33; 
32'd1088: dataIn2 = 32'd22; 
32'd1089: dataIn2 = 32'd27; 
32'd1090: dataIn2 = 32'd63; 
32'd1091: dataIn2 = 32'd59; 
32'd1092: dataIn2 = 32'd31; 
32'd1093: dataIn2 = 32'd4; 
32'd1094: dataIn2 = 32'd98; 
32'd1095: dataIn2 = 32'd37; 
32'd1096: dataIn2 = 32'd16; 
32'd1097: dataIn2 = 32'd84; 
32'd1098: dataIn2 = 32'd26; 
32'd1099: dataIn2 = 32'd80; 
32'd1100: dataIn2 = 32'd50; 
32'd1101: dataIn2 = 32'd23; 
32'd1102: dataIn2 = 32'd43; 
32'd1103: dataIn2 = 32'd2; 
32'd1104: dataIn2 = 32'd46; 
32'd1105: dataIn2 = 32'd26; 
32'd1106: dataIn2 = 32'd31; 
32'd1107: dataIn2 = 32'd32; 
32'd1108: dataIn2 = 32'd6; 
32'd1109: dataIn2 = 32'd41; 
32'd1110: dataIn2 = 32'd47; 
32'd1111: dataIn2 = 32'd69; 
32'd1112: dataIn2 = 32'd0; 
32'd1113: dataIn2 = 32'd39; 
32'd1114: dataIn2 = 32'd4; 
32'd1115: dataIn2 = 32'd59; 
32'd1116: dataIn2 = 32'd45; 
32'd1117: dataIn2 = 32'd0; 
32'd1118: dataIn2 = 32'd57; 
32'd1119: dataIn2 = 32'd48; 
32'd1120: dataIn2 = 32'd85; 
32'd1121: dataIn2 = 32'd97; 
32'd1122: dataIn2 = 32'd48; 
32'd1123: dataIn2 = 32'd100; 
32'd1124: dataIn2 = 32'd14; 
32'd1125: dataIn2 = 32'd23; 
32'd1126: dataIn2 = 32'd90; 
32'd1127: dataIn2 = 32'd4; 
32'd1128: dataIn2 = 32'd35; 
32'd1129: dataIn2 = 32'd85; 
32'd1130: dataIn2 = 32'd6; 
32'd1131: dataIn2 = 32'd87; 
32'd1132: dataIn2 = 32'd16; 
32'd1133: dataIn2 = 32'd74; 
32'd1134: dataIn2 = 32'd10; 
32'd1135: dataIn2 = 32'd57; 
32'd1136: dataIn2 = 32'd61; 
32'd1137: dataIn2 = 32'd1; 
32'd1138: dataIn2 = 32'd36; 
32'd1139: dataIn2 = 32'd100; 
32'd1140: dataIn2 = 32'd1; 
32'd1141: dataIn2 = 32'd41; 
32'd1142: dataIn2 = 32'd59; 
32'd1143: dataIn2 = 32'd14; 
32'd1144: dataIn2 = 32'd66; 
32'd1145: dataIn2 = 32'd47; 
32'd1146: dataIn2 = 32'd100; 
32'd1147: dataIn2 = 32'd85; 
32'd1148: dataIn2 = 32'd32; 
32'd1149: dataIn2 = 32'd1; 
32'd1150: dataIn2 = 32'd4; 
32'd1151: dataIn2 = 32'd33; 
32'd1152: dataIn2 = 32'd88; 
32'd1153: dataIn2 = 32'd64; 
32'd1154: dataIn2 = 32'd21; 
32'd1155: dataIn2 = 32'd24; 
32'd1156: dataIn2 = 32'd48; 
32'd1157: dataIn2 = 32'd44; 
32'd1158: dataIn2 = 32'd61; 
32'd1159: dataIn2 = 32'd95; 
32'd1160: dataIn2 = 32'd9; 
32'd1161: dataIn2 = 32'd22; 
32'd1162: dataIn2 = 32'd100; 
32'd1163: dataIn2 = 32'd15; 
32'd1164: dataIn2 = 32'd58; 
32'd1165: dataIn2 = 32'd43; 
32'd1166: dataIn2 = 32'd17; 
32'd1167: dataIn2 = 32'd5; 
32'd1168: dataIn2 = 32'd71; 
32'd1169: dataIn2 = 32'd66; 
32'd1170: dataIn2 = 32'd66; 
32'd1171: dataIn2 = 32'd83; 
32'd1172: dataIn2 = 32'd19; 
32'd1173: dataIn2 = 32'd95; 
32'd1174: dataIn2 = 32'd45; 
32'd1175: dataIn2 = 32'd100; 
32'd1176: dataIn2 = 32'd8; 
32'd1177: dataIn2 = 32'd28; 
32'd1178: dataIn2 = 32'd91; 
32'd1179: dataIn2 = 32'd6; 
32'd1180: dataIn2 = 32'd22; 
32'd1181: dataIn2 = 32'd66; 
32'd1182: dataIn2 = 32'd85; 
32'd1183: dataIn2 = 32'd8; 
32'd1184: dataIn2 = 32'd42; 
32'd1185: dataIn2 = 32'd31; 
32'd1186: dataIn2 = 32'd28; 
32'd1187: dataIn2 = 32'd73; 
32'd1188: dataIn2 = 32'd100; 
32'd1189: dataIn2 = 32'd4; 
32'd1190: dataIn2 = 32'd93; 
32'd1191: dataIn2 = 32'd79; 
32'd1192: dataIn2 = 32'd29; 
32'd1193: dataIn2 = 32'd14; 
32'd1194: dataIn2 = 32'd30; 
32'd1195: dataIn2 = 32'd12; 
32'd1196: dataIn2 = 32'd95; 
32'd1197: dataIn2 = 32'd17; 
32'd1198: dataIn2 = 32'd94; 
32'd1199: dataIn2 = 32'd48; 
32'd1200: dataIn2 = 32'd99; 
32'd1201: dataIn2 = 32'd71; 
32'd1202: dataIn2 = 32'd29; 
32'd1203: dataIn2 = 32'd85; 
32'd1204: dataIn2 = 32'd38; 
32'd1205: dataIn2 = 32'd10; 
32'd1206: dataIn2 = 32'd80; 
32'd1207: dataIn2 = 32'd34; 
32'd1208: dataIn2 = 32'd10; 
32'd1209: dataIn2 = 32'd97; 
32'd1210: dataIn2 = 32'd61; 
32'd1211: dataIn2 = 32'd96; 
32'd1212: dataIn2 = 32'd19; 
32'd1213: dataIn2 = 32'd96; 
32'd1214: dataIn2 = 32'd0; 
32'd1215: dataIn2 = 32'd48; 
32'd1216: dataIn2 = 32'd73; 
32'd1217: dataIn2 = 32'd24; 
32'd1218: dataIn2 = 32'd100; 
32'd1219: dataIn2 = 32'd95; 
32'd1220: dataIn2 = 32'd57; 
32'd1221: dataIn2 = 32'd98; 
32'd1222: dataIn2 = 32'd98; 
32'd1223: dataIn2 = 32'd62; 
32'd1224: dataIn2 = 32'd25; 
32'd1225: dataIn2 = 32'd59; 
32'd1226: dataIn2 = 32'd22; 
32'd1227: dataIn2 = 32'd5; 
32'd1228: dataIn2 = 32'd38; 
32'd1229: dataIn2 = 32'd74; 
32'd1230: dataIn2 = 32'd40; 
32'd1231: dataIn2 = 32'd6; 
32'd1232: dataIn2 = 32'd35; 
32'd1233: dataIn2 = 32'd93; 
32'd1234: dataIn2 = 32'd32; 
32'd1235: dataIn2 = 32'd27; 
32'd1236: dataIn2 = 32'd8; 
32'd1237: dataIn2 = 32'd41; 
32'd1238: dataIn2 = 32'd11; 
32'd1239: dataIn2 = 32'd100; 
32'd1240: dataIn2 = 32'd77; 
32'd1241: dataIn2 = 32'd85; 
32'd1242: dataIn2 = 32'd14; 
32'd1243: dataIn2 = 32'd49; 
32'd1244: dataIn2 = 32'd42; 
32'd1245: dataIn2 = 32'd19; 
32'd1246: dataIn2 = 32'd92; 
32'd1247: dataIn2 = 32'd18; 
32'd1248: dataIn2 = 32'd5; 
32'd1249: dataIn2 = 32'd24; 
32'd1250: dataIn2 = 32'd32; 
32'd1251: dataIn2 = 32'd74; 
32'd1252: dataIn2 = 32'd8; 
32'd1253: dataIn2 = 32'd20; 
32'd1254: dataIn2 = 32'd71; 
32'd1255: dataIn2 = 32'd76; 
32'd1256: dataIn2 = 32'd44; 
32'd1257: dataIn2 = 32'd59; 
32'd1258: dataIn2 = 32'd95; 
32'd1259: dataIn2 = 32'd7; 
32'd1260: dataIn2 = 32'd85; 
32'd1261: dataIn2 = 32'd69; 
32'd1262: dataIn2 = 32'd9; 
32'd1263: dataIn2 = 32'd54; 
32'd1264: dataIn2 = 32'd85; 
32'd1265: dataIn2 = 32'd93; 
32'd1266: dataIn2 = 32'd14; 
32'd1267: dataIn2 = 32'd69; 
32'd1268: dataIn2 = 32'd1; 
32'd1269: dataIn2 = 32'd61; 
32'd1270: dataIn2 = 32'd6; 
32'd1271: dataIn2 = 32'd37; 
32'd1272: dataIn2 = 32'd41; 
32'd1273: dataIn2 = 32'd44; 
32'd1274: dataIn2 = 32'd28; 
32'd1275: dataIn2 = 32'd10; 
32'd1276: dataIn2 = 32'd27; 
32'd1277: dataIn2 = 32'd14; 
32'd1278: dataIn2 = 32'd54; 
32'd1279: dataIn2 = 32'd6; 
32'd1280: dataIn2 = 32'd12; 
32'd1281: dataIn2 = 32'd86; 
32'd1282: dataIn2 = 32'd60; 
32'd1283: dataIn2 = 32'd61; 
32'd1284: dataIn2 = 32'd37; 
32'd1285: dataIn2 = 32'd36; 
32'd1286: dataIn2 = 32'd89; 
32'd1287: dataIn2 = 32'd30; 
32'd1288: dataIn2 = 32'd80; 
32'd1289: dataIn2 = 32'd71; 
32'd1290: dataIn2 = 32'd93; 
32'd1291: dataIn2 = 32'd45; 
32'd1292: dataIn2 = 32'd100; 
32'd1293: dataIn2 = 32'd55; 
32'd1294: dataIn2 = 32'd36; 
32'd1295: dataIn2 = 32'd54; 
32'd1296: dataIn2 = 32'd24; 
32'd1297: dataIn2 = 32'd31; 
32'd1298: dataIn2 = 32'd29; 
32'd1299: dataIn2 = 32'd76; 
32'd1300: dataIn2 = 32'd17; 
32'd1301: dataIn2 = 32'd18; 
32'd1302: dataIn2 = 32'd2; 
32'd1303: dataIn2 = 32'd81; 
32'd1304: dataIn2 = 32'd65; 
32'd1305: dataIn2 = 32'd6; 
32'd1306: dataIn2 = 32'd58; 
32'd1307: dataIn2 = 32'd5; 
32'd1308: dataIn2 = 32'd31; 
32'd1309: dataIn2 = 32'd39; 
32'd1310: dataIn2 = 32'd44; 
32'd1311: dataIn2 = 32'd71; 
32'd1312: dataIn2 = 32'd59; 
32'd1313: dataIn2 = 32'd60; 
32'd1314: dataIn2 = 32'd38; 
32'd1315: dataIn2 = 32'd51; 
32'd1316: dataIn2 = 32'd56; 
32'd1317: dataIn2 = 32'd69; 
32'd1318: dataIn2 = 32'd57; 
32'd1319: dataIn2 = 32'd36; 
32'd1320: dataIn2 = 32'd12; 
32'd1321: dataIn2 = 32'd38; 
32'd1322: dataIn2 = 32'd25; 
32'd1323: dataIn2 = 32'd77; 
32'd1324: dataIn2 = 32'd78; 
32'd1325: dataIn2 = 32'd8; 
32'd1326: dataIn2 = 32'd33; 
32'd1327: dataIn2 = 32'd100; 
32'd1328: dataIn2 = 32'd21; 
32'd1329: dataIn2 = 32'd69; 
32'd1330: dataIn2 = 32'd24; 
32'd1331: dataIn2 = 32'd10; 
32'd1332: dataIn2 = 32'd96; 
32'd1333: dataIn2 = 32'd43; 
32'd1334: dataIn2 = 32'd10; 
32'd1335: dataIn2 = 32'd50; 
32'd1336: dataIn2 = 32'd68; 
32'd1337: dataIn2 = 32'd60; 
32'd1338: dataIn2 = 32'd24; 
32'd1339: dataIn2 = 32'd67; 
32'd1340: dataIn2 = 32'd71; 
32'd1341: dataIn2 = 32'd72; 
32'd1342: dataIn2 = 32'd87; 
32'd1343: dataIn2 = 32'd5; 
32'd1344: dataIn2 = 32'd46; 
32'd1345: dataIn2 = 32'd45; 
32'd1346: dataIn2 = 32'd25; 
32'd1347: dataIn2 = 32'd50; 
32'd1348: dataIn2 = 32'd91; 
32'd1349: dataIn2 = 32'd2; 
32'd1350: dataIn2 = 32'd55; 
32'd1351: dataIn2 = 32'd76; 
32'd1352: dataIn2 = 32'd30; 
32'd1353: dataIn2 = 32'd99; 
32'd1354: dataIn2 = 32'd4; 
32'd1355: dataIn2 = 32'd42; 
32'd1356: dataIn2 = 32'd48; 
32'd1357: dataIn2 = 32'd95; 
32'd1358: dataIn2 = 32'd74; 
32'd1359: dataIn2 = 32'd68; 
32'd1360: dataIn2 = 32'd20; 
32'd1361: dataIn2 = 32'd30; 
32'd1362: dataIn2 = 32'd72; 
32'd1363: dataIn2 = 32'd43; 
32'd1364: dataIn2 = 32'd3; 
32'd1365: dataIn2 = 32'd67; 
32'd1366: dataIn2 = 32'd56; 
32'd1367: dataIn2 = 32'd71; 
32'd1368: dataIn2 = 32'd78; 
32'd1369: dataIn2 = 32'd72; 
32'd1370: dataIn2 = 32'd33; 
32'd1371: dataIn2 = 32'd1; 
32'd1372: dataIn2 = 32'd31; 
32'd1373: dataIn2 = 32'd26; 
32'd1374: dataIn2 = 32'd47; 
32'd1375: dataIn2 = 32'd78; 
32'd1376: dataIn2 = 32'd69; 
32'd1377: dataIn2 = 32'd33; 
32'd1378: dataIn2 = 32'd49; 
32'd1379: dataIn2 = 32'd54; 
32'd1380: dataIn2 = 32'd28; 
32'd1381: dataIn2 = 32'd0; 
32'd1382: dataIn2 = 32'd87; 
32'd1383: dataIn2 = 32'd38; 
32'd1384: dataIn2 = 32'd95; 
32'd1385: dataIn2 = 32'd26; 
32'd1386: dataIn2 = 32'd25; 
32'd1387: dataIn2 = 32'd73; 
32'd1388: dataIn2 = 32'd1; 
32'd1389: dataIn2 = 32'd1; 
32'd1390: dataIn2 = 32'd75; 
32'd1391: dataIn2 = 32'd100; 
32'd1392: dataIn2 = 32'd33; 
32'd1393: dataIn2 = 32'd22; 
32'd1394: dataIn2 = 32'd31; 
32'd1395: dataIn2 = 32'd74; 
32'd1396: dataIn2 = 32'd41; 
32'd1397: dataIn2 = 32'd22; 
32'd1398: dataIn2 = 32'd82; 
32'd1399: dataIn2 = 32'd75; 
32'd1400: dataIn2 = 32'd0; 
32'd1401: dataIn2 = 32'd6; 
32'd1402: dataIn2 = 32'd20; 
32'd1403: dataIn2 = 32'd68; 
32'd1404: dataIn2 = 32'd12; 
32'd1405: dataIn2 = 32'd41; 
32'd1406: dataIn2 = 32'd94; 
32'd1407: dataIn2 = 32'd18; 
32'd1408: dataIn2 = 32'd43; 
32'd1409: dataIn2 = 32'd52; 
32'd1410: dataIn2 = 32'd47; 
32'd1411: dataIn2 = 32'd23; 
32'd1412: dataIn2 = 32'd32; 
32'd1413: dataIn2 = 32'd91; 
32'd1414: dataIn2 = 32'd6; 
32'd1415: dataIn2 = 32'd45; 
32'd1416: dataIn2 = 32'd67; 
32'd1417: dataIn2 = 32'd38; 
32'd1418: dataIn2 = 32'd83; 
32'd1419: dataIn2 = 32'd78; 
32'd1420: dataIn2 = 32'd21; 
32'd1421: dataIn2 = 32'd73; 
32'd1422: dataIn2 = 32'd80; 
32'd1423: dataIn2 = 32'd97; 
32'd1424: dataIn2 = 32'd91; 
32'd1425: dataIn2 = 32'd87; 
32'd1426: dataIn2 = 32'd16; 
32'd1427: dataIn2 = 32'd45; 
32'd1428: dataIn2 = 32'd79; 
32'd1429: dataIn2 = 32'd89; 
32'd1430: dataIn2 = 32'd21; 
32'd1431: dataIn2 = 32'd2; 
32'd1432: dataIn2 = 32'd61; 
32'd1433: dataIn2 = 32'd5; 
32'd1434: dataIn2 = 32'd60; 
32'd1435: dataIn2 = 32'd12; 
32'd1436: dataIn2 = 32'd79; 
32'd1437: dataIn2 = 32'd66; 
32'd1438: dataIn2 = 32'd67; 
32'd1439: dataIn2 = 32'd86; 
32'd1440: dataIn2 = 32'd12; 
32'd1441: dataIn2 = 32'd53; 
32'd1442: dataIn2 = 32'd12; 
32'd1443: dataIn2 = 32'd94; 
32'd1444: dataIn2 = 32'd20; 
32'd1445: dataIn2 = 32'd51; 
32'd1446: dataIn2 = 32'd61; 
32'd1447: dataIn2 = 32'd88; 
32'd1448: dataIn2 = 32'd27; 
32'd1449: dataIn2 = 32'd23; 
32'd1450: dataIn2 = 32'd31; 
32'd1451: dataIn2 = 32'd4; 
32'd1452: dataIn2 = 32'd68; 
32'd1453: dataIn2 = 32'd72; 
32'd1454: dataIn2 = 32'd14; 
32'd1455: dataIn2 = 32'd38; 
32'd1456: dataIn2 = 32'd33; 
32'd1457: dataIn2 = 32'd60; 
32'd1458: dataIn2 = 32'd11; 
32'd1459: dataIn2 = 32'd2; 
32'd1460: dataIn2 = 32'd36; 
32'd1461: dataIn2 = 32'd67; 
32'd1462: dataIn2 = 32'd11; 
32'd1463: dataIn2 = 32'd90; 
32'd1464: dataIn2 = 32'd51; 
32'd1465: dataIn2 = 32'd32; 
32'd1466: dataIn2 = 32'd31; 
32'd1467: dataIn2 = 32'd13; 
32'd1468: dataIn2 = 32'd19; 
32'd1469: dataIn2 = 32'd91; 
32'd1470: dataIn2 = 32'd1; 
32'd1471: dataIn2 = 32'd43; 
32'd1472: dataIn2 = 32'd19; 
32'd1473: dataIn2 = 32'd54; 
32'd1474: dataIn2 = 32'd26; 
32'd1475: dataIn2 = 32'd53; 
32'd1476: dataIn2 = 32'd45; 
32'd1477: dataIn2 = 32'd95; 
32'd1478: dataIn2 = 32'd16; 
32'd1479: dataIn2 = 32'd50; 
32'd1480: dataIn2 = 32'd6; 
32'd1481: dataIn2 = 32'd88; 
32'd1482: dataIn2 = 32'd62; 
32'd1483: dataIn2 = 32'd3; 
32'd1484: dataIn2 = 32'd51; 
32'd1485: dataIn2 = 32'd28; 
32'd1486: dataIn2 = 32'd59; 
32'd1487: dataIn2 = 32'd84; 
32'd1488: dataIn2 = 32'd39; 
32'd1489: dataIn2 = 32'd8; 
32'd1490: dataIn2 = 32'd72; 
32'd1491: dataIn2 = 32'd56; 
32'd1492: dataIn2 = 32'd44; 
32'd1493: dataIn2 = 32'd36; 
32'd1494: dataIn2 = 32'd29; 
32'd1495: dataIn2 = 32'd29; 
32'd1496: dataIn2 = 32'd66; 
32'd1497: dataIn2 = 32'd90; 
32'd1498: dataIn2 = 32'd52; 
32'd1499: dataIn2 = 32'd62; 
32'd1500: dataIn2 = 32'd97; 
32'd1501: dataIn2 = 32'd1; 
32'd1502: dataIn2 = 32'd83; 
32'd1503: dataIn2 = 32'd46; 
32'd1504: dataIn2 = 32'd11; 
32'd1505: dataIn2 = 32'd13; 
32'd1506: dataIn2 = 32'd92; 
32'd1507: dataIn2 = 32'd46; 
32'd1508: dataIn2 = 32'd51; 
32'd1509: dataIn2 = 32'd95; 
32'd1510: dataIn2 = 32'd100; 
32'd1511: dataIn2 = 32'd66; 
32'd1512: dataIn2 = 32'd1; 
32'd1513: dataIn2 = 32'd97; 
32'd1514: dataIn2 = 32'd84; 
32'd1515: dataIn2 = 32'd52; 
32'd1516: dataIn2 = 32'd98; 
32'd1517: dataIn2 = 32'd31; 
32'd1518: dataIn2 = 32'd77; 
32'd1519: dataIn2 = 32'd26; 
32'd1520: dataIn2 = 32'd33; 
32'd1521: dataIn2 = 32'd27; 
32'd1522: dataIn2 = 32'd24; 
32'd1523: dataIn2 = 32'd67; 
32'd1524: dataIn2 = 32'd35; 
32'd1525: dataIn2 = 32'd75; 
32'd1526: dataIn2 = 32'd43; 
32'd1527: dataIn2 = 32'd81; 
32'd1528: dataIn2 = 32'd44; 
32'd1529: dataIn2 = 32'd2; 
32'd1530: dataIn2 = 32'd37; 
32'd1531: dataIn2 = 32'd22; 
32'd1532: dataIn2 = 32'd41; 
32'd1533: dataIn2 = 32'd62; 
32'd1534: dataIn2 = 32'd53; 
32'd1535: dataIn2 = 32'd23; 
32'd1536: dataIn2 = 32'd97; 
32'd1537: dataIn2 = 32'd19; 
32'd1538: dataIn2 = 32'd51; 
32'd1539: dataIn2 = 32'd88; 
32'd1540: dataIn2 = 32'd53; 
32'd1541: dataIn2 = 32'd10; 
32'd1542: dataIn2 = 32'd56; 
32'd1543: dataIn2 = 32'd76; 
32'd1544: dataIn2 = 32'd49; 
32'd1545: dataIn2 = 32'd27; 
32'd1546: dataIn2 = 32'd38; 
32'd1547: dataIn2 = 32'd99; 
32'd1548: dataIn2 = 32'd16; 
32'd1549: dataIn2 = 32'd87; 
32'd1550: dataIn2 = 32'd26; 
32'd1551: dataIn2 = 32'd26; 
32'd1552: dataIn2 = 32'd32; 
32'd1553: dataIn2 = 32'd51; 
32'd1554: dataIn2 = 32'd2; 
32'd1555: dataIn2 = 32'd47; 
32'd1556: dataIn2 = 32'd5; 
32'd1557: dataIn2 = 32'd18; 
32'd1558: dataIn2 = 32'd52; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_64_70.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
