//32x32 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 717 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd170 ; 
  wdata_col_base = 32'd8870 ; 
  row_base = 32'd95870 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #14520; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd95870: dataIn1 = 32'd0
; 
32'd95871: dataIn1 = 32'd23
; 
32'd95872: dataIn1 = 32'd50
; 
32'd95873: dataIn1 = 32'd70
; 
32'd95874: dataIn1 = 32'd85
; 
32'd95875: dataIn1 = 32'd104
; 
32'd95876: dataIn1 = 32'd126
; 
32'd95877: dataIn1 = 32'd151
; 
32'd95878: dataIn1 = 32'd174
; 
32'd95879: dataIn1 = 32'd200
; 
32'd95880: dataIn1 = 32'd221
; 
32'd95881: dataIn1 = 32'd247
; 
32'd95882: dataIn1 = 32'd269
; 
32'd95883: dataIn1 = 32'd292
; 
32'd95884: dataIn1 = 32'd311
; 
32'd95885: dataIn1 = 32'd334
; 
32'd95886: dataIn1 = 32'd360
; 
32'd95887: dataIn1 = 32'd377
; 
32'd95888: dataIn1 = 32'd395
; 
32'd95889: dataIn1 = 32'd414
; 
32'd95890: dataIn1 = 32'd437
; 
32'd95891: dataIn1 = 32'd462
; 
32'd95892: dataIn1 = 32'd483
; 
32'd95893: dataIn1 = 32'd507
; 
32'd95894: dataIn1 = 32'd527
; 
32'd95895: dataIn1 = 32'd549
; 
32'd95896: dataIn1 = 32'd573
; 
32'd95897: dataIn1 = 32'd593
; 
32'd95898: dataIn1 = 32'd615
; 
32'd95899: dataIn1 = 32'd633
; 
32'd95900: dataIn1 = 32'd658
; 
32'd95901: dataIn1 = 32'd680
; 
32'd95902: dataIn1 = 32'd699
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd8870: dataIn1 = 32'd0
; 
32'd8871: dataIn1 = 32'd23
; 
32'd8872: dataIn1 = 32'd50
; 
32'd8873: dataIn1 = 32'd70
; 
32'd8874: dataIn1 = 32'd85
; 
32'd8875: dataIn1 = 32'd104
; 
32'd8876: dataIn1 = 32'd126
; 
32'd8877: dataIn1 = 32'd151
; 
32'd8878: dataIn1 = 32'd174
; 
32'd8879: dataIn1 = 32'd200
; 
32'd8880: dataIn1 = 32'd221
; 
32'd8881: dataIn1 = 32'd247
; 
32'd8882: dataIn1 = 32'd269
; 
32'd8883: dataIn1 = 32'd292
; 
32'd8884: dataIn1 = 32'd311
; 
32'd8885: dataIn1 = 32'd334
; 
32'd8886: dataIn1 = 32'd360
; 
32'd8887: dataIn1 = 32'd377
; 
32'd8888: dataIn1 = 32'd395
; 
32'd8889: dataIn1 = 32'd414
; 
32'd8890: dataIn1 = 32'd437
; 
32'd8891: dataIn1 = 32'd462
; 
32'd8892: dataIn1 = 32'd483
; 
32'd8893: dataIn1 = 32'd507
; 
32'd8894: dataIn1 = 32'd527
; 
32'd8895: dataIn1 = 32'd549
; 
32'd8896: dataIn1 = 32'd573
; 
32'd8897: dataIn1 = 32'd593
; 
32'd8898: dataIn1 = 32'd615
; 
32'd8899: dataIn1 = 32'd633
; 
32'd8900: dataIn1 = 32'd658
; 
32'd8901: dataIn1 = 32'd680
; 
32'd8902: dataIn1 = 32'd699
; 
32'd8903: dataIn1 = 32'd0
; 
32'd8904: dataIn1 = 32'd1
; 
32'd8905: dataIn1 = 32'd2
; 
32'd8906: dataIn1 = 32'd3
; 
32'd8907: dataIn1 = 32'd5
; 
32'd8908: dataIn1 = 32'd6
; 
32'd8909: dataIn1 = 32'd8
; 
32'd8910: dataIn1 = 32'd9
; 
32'd8911: dataIn1 = 32'd10
; 
32'd8912: dataIn1 = 32'd12
; 
32'd8913: dataIn1 = 32'd13
; 
32'd8914: dataIn1 = 32'd14
; 
32'd8915: dataIn1 = 32'd16
; 
32'd8916: dataIn1 = 32'd17
; 
32'd8917: dataIn1 = 32'd18
; 
32'd8918: dataIn1 = 32'd19
; 
32'd8919: dataIn1 = 32'd20
; 
32'd8920: dataIn1 = 32'd21
; 
32'd8921: dataIn1 = 32'd22
; 
32'd8922: dataIn1 = 32'd24
; 
32'd8923: dataIn1 = 32'd26
; 
32'd8924: dataIn1 = 32'd27
; 
32'd8925: dataIn1 = 32'd28
; 
32'd8926: dataIn1 = 32'd0
; 
32'd8927: dataIn1 = 32'd1
; 
32'd8928: dataIn1 = 32'd2
; 
32'd8929: dataIn1 = 32'd3
; 
32'd8930: dataIn1 = 32'd6
; 
32'd8931: dataIn1 = 32'd7
; 
32'd8932: dataIn1 = 32'd8
; 
32'd8933: dataIn1 = 32'd9
; 
32'd8934: dataIn1 = 32'd10
; 
32'd8935: dataIn1 = 32'd12
; 
32'd8936: dataIn1 = 32'd13
; 
32'd8937: dataIn1 = 32'd14
; 
32'd8938: dataIn1 = 32'd15
; 
32'd8939: dataIn1 = 32'd16
; 
32'd8940: dataIn1 = 32'd17
; 
32'd8941: dataIn1 = 32'd18
; 
32'd8942: dataIn1 = 32'd19
; 
32'd8943: dataIn1 = 32'd21
; 
32'd8944: dataIn1 = 32'd22
; 
32'd8945: dataIn1 = 32'd23
; 
32'd8946: dataIn1 = 32'd24
; 
32'd8947: dataIn1 = 32'd25
; 
32'd8948: dataIn1 = 32'd26
; 
32'd8949: dataIn1 = 32'd27
; 
32'd8950: dataIn1 = 32'd29
; 
32'd8951: dataIn1 = 32'd30
; 
32'd8952: dataIn1 = 32'd31
; 
32'd8953: dataIn1 = 32'd0
; 
32'd8954: dataIn1 = 32'd3
; 
32'd8955: dataIn1 = 32'd4
; 
32'd8956: dataIn1 = 32'd6
; 
32'd8957: dataIn1 = 32'd7
; 
32'd8958: dataIn1 = 32'd9
; 
32'd8959: dataIn1 = 32'd11
; 
32'd8960: dataIn1 = 32'd12
; 
32'd8961: dataIn1 = 32'd13
; 
32'd8962: dataIn1 = 32'd15
; 
32'd8963: dataIn1 = 32'd17
; 
32'd8964: dataIn1 = 32'd19
; 
32'd8965: dataIn1 = 32'd20
; 
32'd8966: dataIn1 = 32'd22
; 
32'd8967: dataIn1 = 32'd23
; 
32'd8968: dataIn1 = 32'd24
; 
32'd8969: dataIn1 = 32'd25
; 
32'd8970: dataIn1 = 32'd26
; 
32'd8971: dataIn1 = 32'd27
; 
32'd8972: dataIn1 = 32'd30
; 
32'd8973: dataIn1 = 32'd0
; 
32'd8974: dataIn1 = 32'd2
; 
32'd8975: dataIn1 = 32'd5
; 
32'd8976: dataIn1 = 32'd6
; 
32'd8977: dataIn1 = 32'd8
; 
32'd8978: dataIn1 = 32'd9
; 
32'd8979: dataIn1 = 32'd11
; 
32'd8980: dataIn1 = 32'd14
; 
32'd8981: dataIn1 = 32'd15
; 
32'd8982: dataIn1 = 32'd17
; 
32'd8983: dataIn1 = 32'd18
; 
32'd8984: dataIn1 = 32'd22
; 
32'd8985: dataIn1 = 32'd23
; 
32'd8986: dataIn1 = 32'd25
; 
32'd8987: dataIn1 = 32'd27
; 
32'd8988: dataIn1 = 32'd0
; 
32'd8989: dataIn1 = 32'd1
; 
32'd8990: dataIn1 = 32'd5
; 
32'd8991: dataIn1 = 32'd7
; 
32'd8992: dataIn1 = 32'd8
; 
32'd8993: dataIn1 = 32'd9
; 
32'd8994: dataIn1 = 32'd10
; 
32'd8995: dataIn1 = 32'd11
; 
32'd8996: dataIn1 = 32'd12
; 
32'd8997: dataIn1 = 32'd13
; 
32'd8998: dataIn1 = 32'd14
; 
32'd8999: dataIn1 = 32'd22
; 
32'd9000: dataIn1 = 32'd23
; 
32'd9001: dataIn1 = 32'd24
; 
32'd9002: dataIn1 = 32'd25
; 
32'd9003: dataIn1 = 32'd26
; 
32'd9004: dataIn1 = 32'd28
; 
32'd9005: dataIn1 = 32'd29
; 
32'd9006: dataIn1 = 32'd31
; 
32'd9007: dataIn1 = 32'd2
; 
32'd9008: dataIn1 = 32'd3
; 
32'd9009: dataIn1 = 32'd4
; 
32'd9010: dataIn1 = 32'd7
; 
32'd9011: dataIn1 = 32'd8
; 
32'd9012: dataIn1 = 32'd9
; 
32'd9013: dataIn1 = 32'd10
; 
32'd9014: dataIn1 = 32'd12
; 
32'd9015: dataIn1 = 32'd13
; 
32'd9016: dataIn1 = 32'd14
; 
32'd9017: dataIn1 = 32'd16
; 
32'd9018: dataIn1 = 32'd17
; 
32'd9019: dataIn1 = 32'd19
; 
32'd9020: dataIn1 = 32'd20
; 
32'd9021: dataIn1 = 32'd21
; 
32'd9022: dataIn1 = 32'd22
; 
32'd9023: dataIn1 = 32'd23
; 
32'd9024: dataIn1 = 32'd25
; 
32'd9025: dataIn1 = 32'd26
; 
32'd9026: dataIn1 = 32'd27
; 
32'd9027: dataIn1 = 32'd29
; 
32'd9028: dataIn1 = 32'd31
; 
32'd9029: dataIn1 = 32'd0
; 
32'd9030: dataIn1 = 32'd1
; 
32'd9031: dataIn1 = 32'd2
; 
32'd9032: dataIn1 = 32'd3
; 
32'd9033: dataIn1 = 32'd4
; 
32'd9034: dataIn1 = 32'd5
; 
32'd9035: dataIn1 = 32'd9
; 
32'd9036: dataIn1 = 32'd10
; 
32'd9037: dataIn1 = 32'd11
; 
32'd9038: dataIn1 = 32'd12
; 
32'd9039: dataIn1 = 32'd13
; 
32'd9040: dataIn1 = 32'd14
; 
32'd9041: dataIn1 = 32'd15
; 
32'd9042: dataIn1 = 32'd16
; 
32'd9043: dataIn1 = 32'd17
; 
32'd9044: dataIn1 = 32'd19
; 
32'd9045: dataIn1 = 32'd20
; 
32'd9046: dataIn1 = 32'd22
; 
32'd9047: dataIn1 = 32'd23
; 
32'd9048: dataIn1 = 32'd25
; 
32'd9049: dataIn1 = 32'd26
; 
32'd9050: dataIn1 = 32'd27
; 
32'd9051: dataIn1 = 32'd28
; 
32'd9052: dataIn1 = 32'd29
; 
32'd9053: dataIn1 = 32'd30
; 
32'd9054: dataIn1 = 32'd0
; 
32'd9055: dataIn1 = 32'd1
; 
32'd9056: dataIn1 = 32'd2
; 
32'd9057: dataIn1 = 32'd4
; 
32'd9058: dataIn1 = 32'd5
; 
32'd9059: dataIn1 = 32'd6
; 
32'd9060: dataIn1 = 32'd7
; 
32'd9061: dataIn1 = 32'd8
; 
32'd9062: dataIn1 = 32'd9
; 
32'd9063: dataIn1 = 32'd11
; 
32'd9064: dataIn1 = 32'd12
; 
32'd9065: dataIn1 = 32'd13
; 
32'd9066: dataIn1 = 32'd14
; 
32'd9067: dataIn1 = 32'd15
; 
32'd9068: dataIn1 = 32'd16
; 
32'd9069: dataIn1 = 32'd17
; 
32'd9070: dataIn1 = 32'd20
; 
32'd9071: dataIn1 = 32'd21
; 
32'd9072: dataIn1 = 32'd22
; 
32'd9073: dataIn1 = 32'd25
; 
32'd9074: dataIn1 = 32'd26
; 
32'd9075: dataIn1 = 32'd28
; 
32'd9076: dataIn1 = 32'd29
; 
32'd9077: dataIn1 = 32'd0
; 
32'd9078: dataIn1 = 32'd1
; 
32'd9079: dataIn1 = 32'd2
; 
32'd9080: dataIn1 = 32'd4
; 
32'd9081: dataIn1 = 32'd5
; 
32'd9082: dataIn1 = 32'd6
; 
32'd9083: dataIn1 = 32'd7
; 
32'd9084: dataIn1 = 32'd8
; 
32'd9085: dataIn1 = 32'd9
; 
32'd9086: dataIn1 = 32'd10
; 
32'd9087: dataIn1 = 32'd12
; 
32'd9088: dataIn1 = 32'd14
; 
32'd9089: dataIn1 = 32'd15
; 
32'd9090: dataIn1 = 32'd16
; 
32'd9091: dataIn1 = 32'd18
; 
32'd9092: dataIn1 = 32'd19
; 
32'd9093: dataIn1 = 32'd20
; 
32'd9094: dataIn1 = 32'd21
; 
32'd9095: dataIn1 = 32'd22
; 
32'd9096: dataIn1 = 32'd23
; 
32'd9097: dataIn1 = 32'd25
; 
32'd9098: dataIn1 = 32'd26
; 
32'd9099: dataIn1 = 32'd27
; 
32'd9100: dataIn1 = 32'd28
; 
32'd9101: dataIn1 = 32'd29
; 
32'd9102: dataIn1 = 32'd30
; 
32'd9103: dataIn1 = 32'd0
; 
32'd9104: dataIn1 = 32'd2
; 
32'd9105: dataIn1 = 32'd3
; 
32'd9106: dataIn1 = 32'd4
; 
32'd9107: dataIn1 = 32'd5
; 
32'd9108: dataIn1 = 32'd6
; 
32'd9109: dataIn1 = 32'd8
; 
32'd9110: dataIn1 = 32'd9
; 
32'd9111: dataIn1 = 32'd10
; 
32'd9112: dataIn1 = 32'd11
; 
32'd9113: dataIn1 = 32'd12
; 
32'd9114: dataIn1 = 32'd15
; 
32'd9115: dataIn1 = 32'd17
; 
32'd9116: dataIn1 = 32'd18
; 
32'd9117: dataIn1 = 32'd19
; 
32'd9118: dataIn1 = 32'd22
; 
32'd9119: dataIn1 = 32'd26
; 
32'd9120: dataIn1 = 32'd27
; 
32'd9121: dataIn1 = 32'd28
; 
32'd9122: dataIn1 = 32'd29
; 
32'd9123: dataIn1 = 32'd31
; 
32'd9124: dataIn1 = 32'd0
; 
32'd9125: dataIn1 = 32'd1
; 
32'd9126: dataIn1 = 32'd2
; 
32'd9127: dataIn1 = 32'd4
; 
32'd9128: dataIn1 = 32'd5
; 
32'd9129: dataIn1 = 32'd6
; 
32'd9130: dataIn1 = 32'd7
; 
32'd9131: dataIn1 = 32'd11
; 
32'd9132: dataIn1 = 32'd12
; 
32'd9133: dataIn1 = 32'd13
; 
32'd9134: dataIn1 = 32'd14
; 
32'd9135: dataIn1 = 32'd15
; 
32'd9136: dataIn1 = 32'd16
; 
32'd9137: dataIn1 = 32'd17
; 
32'd9138: dataIn1 = 32'd18
; 
32'd9139: dataIn1 = 32'd19
; 
32'd9140: dataIn1 = 32'd21
; 
32'd9141: dataIn1 = 32'd22
; 
32'd9142: dataIn1 = 32'd23
; 
32'd9143: dataIn1 = 32'd24
; 
32'd9144: dataIn1 = 32'd25
; 
32'd9145: dataIn1 = 32'd26
; 
32'd9146: dataIn1 = 32'd27
; 
32'd9147: dataIn1 = 32'd29
; 
32'd9148: dataIn1 = 32'd30
; 
32'd9149: dataIn1 = 32'd31
; 
32'd9150: dataIn1 = 32'd0
; 
32'd9151: dataIn1 = 32'd1
; 
32'd9152: dataIn1 = 32'd2
; 
32'd9153: dataIn1 = 32'd3
; 
32'd9154: dataIn1 = 32'd4
; 
32'd9155: dataIn1 = 32'd5
; 
32'd9156: dataIn1 = 32'd6
; 
32'd9157: dataIn1 = 32'd8
; 
32'd9158: dataIn1 = 32'd10
; 
32'd9159: dataIn1 = 32'd11
; 
32'd9160: dataIn1 = 32'd12
; 
32'd9161: dataIn1 = 32'd13
; 
32'd9162: dataIn1 = 32'd15
; 
32'd9163: dataIn1 = 32'd16
; 
32'd9164: dataIn1 = 32'd19
; 
32'd9165: dataIn1 = 32'd20
; 
32'd9166: dataIn1 = 32'd22
; 
32'd9167: dataIn1 = 32'd24
; 
32'd9168: dataIn1 = 32'd27
; 
32'd9169: dataIn1 = 32'd28
; 
32'd9170: dataIn1 = 32'd29
; 
32'd9171: dataIn1 = 32'd30
; 
32'd9172: dataIn1 = 32'd0
; 
32'd9173: dataIn1 = 32'd1
; 
32'd9174: dataIn1 = 32'd2
; 
32'd9175: dataIn1 = 32'd3
; 
32'd9176: dataIn1 = 32'd5
; 
32'd9177: dataIn1 = 32'd6
; 
32'd9178: dataIn1 = 32'd7
; 
32'd9179: dataIn1 = 32'd8
; 
32'd9180: dataIn1 = 32'd9
; 
32'd9181: dataIn1 = 32'd10
; 
32'd9182: dataIn1 = 32'd11
; 
32'd9183: dataIn1 = 32'd12
; 
32'd9184: dataIn1 = 32'd14
; 
32'd9185: dataIn1 = 32'd15
; 
32'd9186: dataIn1 = 32'd17
; 
32'd9187: dataIn1 = 32'd18
; 
32'd9188: dataIn1 = 32'd21
; 
32'd9189: dataIn1 = 32'd26
; 
32'd9190: dataIn1 = 32'd27
; 
32'd9191: dataIn1 = 32'd28
; 
32'd9192: dataIn1 = 32'd29
; 
32'd9193: dataIn1 = 32'd30
; 
32'd9194: dataIn1 = 32'd31
; 
32'd9195: dataIn1 = 32'd1
; 
32'd9196: dataIn1 = 32'd2
; 
32'd9197: dataIn1 = 32'd3
; 
32'd9198: dataIn1 = 32'd4
; 
32'd9199: dataIn1 = 32'd5
; 
32'd9200: dataIn1 = 32'd7
; 
32'd9201: dataIn1 = 32'd11
; 
32'd9202: dataIn1 = 32'd12
; 
32'd9203: dataIn1 = 32'd14
; 
32'd9204: dataIn1 = 32'd16
; 
32'd9205: dataIn1 = 32'd17
; 
32'd9206: dataIn1 = 32'd18
; 
32'd9207: dataIn1 = 32'd22
; 
32'd9208: dataIn1 = 32'd23
; 
32'd9209: dataIn1 = 32'd26
; 
32'd9210: dataIn1 = 32'd27
; 
32'd9211: dataIn1 = 32'd28
; 
32'd9212: dataIn1 = 32'd30
; 
32'd9213: dataIn1 = 32'd31
; 
32'd9214: dataIn1 = 32'd1
; 
32'd9215: dataIn1 = 32'd2
; 
32'd9216: dataIn1 = 32'd3
; 
32'd9217: dataIn1 = 32'd4
; 
32'd9218: dataIn1 = 32'd9
; 
32'd9219: dataIn1 = 32'd10
; 
32'd9220: dataIn1 = 32'd11
; 
32'd9221: dataIn1 = 32'd13
; 
32'd9222: dataIn1 = 32'd14
; 
32'd9223: dataIn1 = 32'd15
; 
32'd9224: dataIn1 = 32'd16
; 
32'd9225: dataIn1 = 32'd17
; 
32'd9226: dataIn1 = 32'd19
; 
32'd9227: dataIn1 = 32'd20
; 
32'd9228: dataIn1 = 32'd21
; 
32'd9229: dataIn1 = 32'd22
; 
32'd9230: dataIn1 = 32'd23
; 
32'd9231: dataIn1 = 32'd24
; 
32'd9232: dataIn1 = 32'd25
; 
32'd9233: dataIn1 = 32'd28
; 
32'd9234: dataIn1 = 32'd29
; 
32'd9235: dataIn1 = 32'd30
; 
32'd9236: dataIn1 = 32'd31
; 
32'd9237: dataIn1 = 32'd0
; 
32'd9238: dataIn1 = 32'd1
; 
32'd9239: dataIn1 = 32'd2
; 
32'd9240: dataIn1 = 32'd3
; 
32'd9241: dataIn1 = 32'd4
; 
32'd9242: dataIn1 = 32'd5
; 
32'd9243: dataIn1 = 32'd6
; 
32'd9244: dataIn1 = 32'd7
; 
32'd9245: dataIn1 = 32'd8
; 
32'd9246: dataIn1 = 32'd10
; 
32'd9247: dataIn1 = 32'd11
; 
32'd9248: dataIn1 = 32'd12
; 
32'd9249: dataIn1 = 32'd14
; 
32'd9250: dataIn1 = 32'd15
; 
32'd9251: dataIn1 = 32'd16
; 
32'd9252: dataIn1 = 32'd17
; 
32'd9253: dataIn1 = 32'd19
; 
32'd9254: dataIn1 = 32'd20
; 
32'd9255: dataIn1 = 32'd21
; 
32'd9256: dataIn1 = 32'd22
; 
32'd9257: dataIn1 = 32'd23
; 
32'd9258: dataIn1 = 32'd25
; 
32'd9259: dataIn1 = 32'd27
; 
32'd9260: dataIn1 = 32'd28
; 
32'd9261: dataIn1 = 32'd30
; 
32'd9262: dataIn1 = 32'd31
; 
32'd9263: dataIn1 = 32'd3
; 
32'd9264: dataIn1 = 32'd4
; 
32'd9265: dataIn1 = 32'd6
; 
32'd9266: dataIn1 = 32'd8
; 
32'd9267: dataIn1 = 32'd9
; 
32'd9268: dataIn1 = 32'd11
; 
32'd9269: dataIn1 = 32'd12
; 
32'd9270: dataIn1 = 32'd15
; 
32'd9271: dataIn1 = 32'd21
; 
32'd9272: dataIn1 = 32'd22
; 
32'd9273: dataIn1 = 32'd23
; 
32'd9274: dataIn1 = 32'd24
; 
32'd9275: dataIn1 = 32'd26
; 
32'd9276: dataIn1 = 32'd27
; 
32'd9277: dataIn1 = 32'd28
; 
32'd9278: dataIn1 = 32'd29
; 
32'd9279: dataIn1 = 32'd30
; 
32'd9280: dataIn1 = 32'd0
; 
32'd9281: dataIn1 = 32'd1
; 
32'd9282: dataIn1 = 32'd5
; 
32'd9283: dataIn1 = 32'd6
; 
32'd9284: dataIn1 = 32'd7
; 
32'd9285: dataIn1 = 32'd8
; 
32'd9286: dataIn1 = 32'd9
; 
32'd9287: dataIn1 = 32'd10
; 
32'd9288: dataIn1 = 32'd11
; 
32'd9289: dataIn1 = 32'd12
; 
32'd9290: dataIn1 = 32'd13
; 
32'd9291: dataIn1 = 32'd16
; 
32'd9292: dataIn1 = 32'd18
; 
32'd9293: dataIn1 = 32'd20
; 
32'd9294: dataIn1 = 32'd22
; 
32'd9295: dataIn1 = 32'd23
; 
32'd9296: dataIn1 = 32'd25
; 
32'd9297: dataIn1 = 32'd26
; 
32'd9298: dataIn1 = 32'd1
; 
32'd9299: dataIn1 = 32'd2
; 
32'd9300: dataIn1 = 32'd4
; 
32'd9301: dataIn1 = 32'd5
; 
32'd9302: dataIn1 = 32'd6
; 
32'd9303: dataIn1 = 32'd10
; 
32'd9304: dataIn1 = 32'd12
; 
32'd9305: dataIn1 = 32'd14
; 
32'd9306: dataIn1 = 32'd15
; 
32'd9307: dataIn1 = 32'd16
; 
32'd9308: dataIn1 = 32'd18
; 
32'd9309: dataIn1 = 32'd19
; 
32'd9310: dataIn1 = 32'd20
; 
32'd9311: dataIn1 = 32'd22
; 
32'd9312: dataIn1 = 32'd24
; 
32'd9313: dataIn1 = 32'd25
; 
32'd9314: dataIn1 = 32'd26
; 
32'd9315: dataIn1 = 32'd29
; 
32'd9316: dataIn1 = 32'd31
; 
32'd9317: dataIn1 = 32'd1
; 
32'd9318: dataIn1 = 32'd2
; 
32'd9319: dataIn1 = 32'd3
; 
32'd9320: dataIn1 = 32'd5
; 
32'd9321: dataIn1 = 32'd6
; 
32'd9322: dataIn1 = 32'd9
; 
32'd9323: dataIn1 = 32'd10
; 
32'd9324: dataIn1 = 32'd11
; 
32'd9325: dataIn1 = 32'd12
; 
32'd9326: dataIn1 = 32'd15
; 
32'd9327: dataIn1 = 32'd16
; 
32'd9328: dataIn1 = 32'd17
; 
32'd9329: dataIn1 = 32'd20
; 
32'd9330: dataIn1 = 32'd21
; 
32'd9331: dataIn1 = 32'd22
; 
32'd9332: dataIn1 = 32'd23
; 
32'd9333: dataIn1 = 32'd24
; 
32'd9334: dataIn1 = 32'd26
; 
32'd9335: dataIn1 = 32'd27
; 
32'd9336: dataIn1 = 32'd28
; 
32'd9337: dataIn1 = 32'd29
; 
32'd9338: dataIn1 = 32'd30
; 
32'd9339: dataIn1 = 32'd31
; 
32'd9340: dataIn1 = 32'd1
; 
32'd9341: dataIn1 = 32'd2
; 
32'd9342: dataIn1 = 32'd3
; 
32'd9343: dataIn1 = 32'd4
; 
32'd9344: dataIn1 = 32'd5
; 
32'd9345: dataIn1 = 32'd8
; 
32'd9346: dataIn1 = 32'd9
; 
32'd9347: dataIn1 = 32'd11
; 
32'd9348: dataIn1 = 32'd13
; 
32'd9349: dataIn1 = 32'd14
; 
32'd9350: dataIn1 = 32'd15
; 
32'd9351: dataIn1 = 32'd17
; 
32'd9352: dataIn1 = 32'd18
; 
32'd9353: dataIn1 = 32'd19
; 
32'd9354: dataIn1 = 32'd21
; 
32'd9355: dataIn1 = 32'd22
; 
32'd9356: dataIn1 = 32'd23
; 
32'd9357: dataIn1 = 32'd24
; 
32'd9358: dataIn1 = 32'd25
; 
32'd9359: dataIn1 = 32'd26
; 
32'd9360: dataIn1 = 32'd27
; 
32'd9361: dataIn1 = 32'd28
; 
32'd9362: dataIn1 = 32'd29
; 
32'd9363: dataIn1 = 32'd30
; 
32'd9364: dataIn1 = 32'd31
; 
32'd9365: dataIn1 = 32'd1
; 
32'd9366: dataIn1 = 32'd2
; 
32'd9367: dataIn1 = 32'd4
; 
32'd9368: dataIn1 = 32'd6
; 
32'd9369: dataIn1 = 32'd7
; 
32'd9370: dataIn1 = 32'd10
; 
32'd9371: dataIn1 = 32'd11
; 
32'd9372: dataIn1 = 32'd12
; 
32'd9373: dataIn1 = 32'd13
; 
32'd9374: dataIn1 = 32'd15
; 
32'd9375: dataIn1 = 32'd17
; 
32'd9376: dataIn1 = 32'd18
; 
32'd9377: dataIn1 = 32'd19
; 
32'd9378: dataIn1 = 32'd20
; 
32'd9379: dataIn1 = 32'd21
; 
32'd9380: dataIn1 = 32'd22
; 
32'd9381: dataIn1 = 32'd23
; 
32'd9382: dataIn1 = 32'd24
; 
32'd9383: dataIn1 = 32'd25
; 
32'd9384: dataIn1 = 32'd28
; 
32'd9385: dataIn1 = 32'd30
; 
32'd9386: dataIn1 = 32'd0
; 
32'd9387: dataIn1 = 32'd2
; 
32'd9388: dataIn1 = 32'd4
; 
32'd9389: dataIn1 = 32'd5
; 
32'd9390: dataIn1 = 32'd6
; 
32'd9391: dataIn1 = 32'd7
; 
32'd9392: dataIn1 = 32'd8
; 
32'd9393: dataIn1 = 32'd9
; 
32'd9394: dataIn1 = 32'd10
; 
32'd9395: dataIn1 = 32'd12
; 
32'd9396: dataIn1 = 32'd13
; 
32'd9397: dataIn1 = 32'd15
; 
32'd9398: dataIn1 = 32'd16
; 
32'd9399: dataIn1 = 32'd17
; 
32'd9400: dataIn1 = 32'd19
; 
32'd9401: dataIn1 = 32'd20
; 
32'd9402: dataIn1 = 32'd21
; 
32'd9403: dataIn1 = 32'd23
; 
32'd9404: dataIn1 = 32'd24
; 
32'd9405: dataIn1 = 32'd25
; 
32'd9406: dataIn1 = 32'd28
; 
32'd9407: dataIn1 = 32'd29
; 
32'd9408: dataIn1 = 32'd30
; 
32'd9409: dataIn1 = 32'd31
; 
32'd9410: dataIn1 = 32'd0
; 
32'd9411: dataIn1 = 32'd1
; 
32'd9412: dataIn1 = 32'd2
; 
32'd9413: dataIn1 = 32'd3
; 
32'd9414: dataIn1 = 32'd8
; 
32'd9415: dataIn1 = 32'd11
; 
32'd9416: dataIn1 = 32'd12
; 
32'd9417: dataIn1 = 32'd13
; 
32'd9418: dataIn1 = 32'd14
; 
32'd9419: dataIn1 = 32'd16
; 
32'd9420: dataIn1 = 32'd17
; 
32'd9421: dataIn1 = 32'd18
; 
32'd9422: dataIn1 = 32'd20
; 
32'd9423: dataIn1 = 32'd21
; 
32'd9424: dataIn1 = 32'd25
; 
32'd9425: dataIn1 = 32'd26
; 
32'd9426: dataIn1 = 32'd28
; 
32'd9427: dataIn1 = 32'd29
; 
32'd9428: dataIn1 = 32'd30
; 
32'd9429: dataIn1 = 32'd31
; 
32'd9430: dataIn1 = 32'd1
; 
32'd9431: dataIn1 = 32'd2
; 
32'd9432: dataIn1 = 32'd3
; 
32'd9433: dataIn1 = 32'd4
; 
32'd9434: dataIn1 = 32'd5
; 
32'd9435: dataIn1 = 32'd6
; 
32'd9436: dataIn1 = 32'd8
; 
32'd9437: dataIn1 = 32'd9
; 
32'd9438: dataIn1 = 32'd10
; 
32'd9439: dataIn1 = 32'd11
; 
32'd9440: dataIn1 = 32'd12
; 
32'd9441: dataIn1 = 32'd13
; 
32'd9442: dataIn1 = 32'd16
; 
32'd9443: dataIn1 = 32'd17
; 
32'd9444: dataIn1 = 32'd18
; 
32'd9445: dataIn1 = 32'd19
; 
32'd9446: dataIn1 = 32'd20
; 
32'd9447: dataIn1 = 32'd23
; 
32'd9448: dataIn1 = 32'd25
; 
32'd9449: dataIn1 = 32'd26
; 
32'd9450: dataIn1 = 32'd29
; 
32'd9451: dataIn1 = 32'd31
; 
32'd9452: dataIn1 = 32'd0
; 
32'd9453: dataIn1 = 32'd1
; 
32'd9454: dataIn1 = 32'd2
; 
32'd9455: dataIn1 = 32'd3
; 
32'd9456: dataIn1 = 32'd6
; 
32'd9457: dataIn1 = 32'd7
; 
32'd9458: dataIn1 = 32'd9
; 
32'd9459: dataIn1 = 32'd10
; 
32'd9460: dataIn1 = 32'd11
; 
32'd9461: dataIn1 = 32'd12
; 
32'd9462: dataIn1 = 32'd14
; 
32'd9463: dataIn1 = 32'd15
; 
32'd9464: dataIn1 = 32'd17
; 
32'd9465: dataIn1 = 32'd19
; 
32'd9466: dataIn1 = 32'd20
; 
32'd9467: dataIn1 = 32'd21
; 
32'd9468: dataIn1 = 32'd22
; 
32'd9469: dataIn1 = 32'd23
; 
32'd9470: dataIn1 = 32'd25
; 
32'd9471: dataIn1 = 32'd26
; 
32'd9472: dataIn1 = 32'd27
; 
32'd9473: dataIn1 = 32'd28
; 
32'd9474: dataIn1 = 32'd29
; 
32'd9475: dataIn1 = 32'd30
; 
32'd9476: dataIn1 = 32'd0
; 
32'd9477: dataIn1 = 32'd2
; 
32'd9478: dataIn1 = 32'd6
; 
32'd9479: dataIn1 = 32'd7
; 
32'd9480: dataIn1 = 32'd8
; 
32'd9481: dataIn1 = 32'd9
; 
32'd9482: dataIn1 = 32'd12
; 
32'd9483: dataIn1 = 32'd13
; 
32'd9484: dataIn1 = 32'd14
; 
32'd9485: dataIn1 = 32'd15
; 
32'd9486: dataIn1 = 32'd16
; 
32'd9487: dataIn1 = 32'd18
; 
32'd9488: dataIn1 = 32'd19
; 
32'd9489: dataIn1 = 32'd20
; 
32'd9490: dataIn1 = 32'd21
; 
32'd9491: dataIn1 = 32'd22
; 
32'd9492: dataIn1 = 32'd25
; 
32'd9493: dataIn1 = 32'd27
; 
32'd9494: dataIn1 = 32'd29
; 
32'd9495: dataIn1 = 32'd30
; 
32'd9496: dataIn1 = 32'd0
; 
32'd9497: dataIn1 = 32'd1
; 
32'd9498: dataIn1 = 32'd2
; 
32'd9499: dataIn1 = 32'd3
; 
32'd9500: dataIn1 = 32'd5
; 
32'd9501: dataIn1 = 32'd9
; 
32'd9502: dataIn1 = 32'd11
; 
32'd9503: dataIn1 = 32'd12
; 
32'd9504: dataIn1 = 32'd14
; 
32'd9505: dataIn1 = 32'd15
; 
32'd9506: dataIn1 = 32'd16
; 
32'd9507: dataIn1 = 32'd17
; 
32'd9508: dataIn1 = 32'd18
; 
32'd9509: dataIn1 = 32'd20
; 
32'd9510: dataIn1 = 32'd22
; 
32'd9511: dataIn1 = 32'd23
; 
32'd9512: dataIn1 = 32'd25
; 
32'd9513: dataIn1 = 32'd27
; 
32'd9514: dataIn1 = 32'd28
; 
32'd9515: dataIn1 = 32'd29
; 
32'd9516: dataIn1 = 32'd30
; 
32'd9517: dataIn1 = 32'd31
; 
32'd9518: dataIn1 = 32'd0
; 
32'd9519: dataIn1 = 32'd1
; 
32'd9520: dataIn1 = 32'd3
; 
32'd9521: dataIn1 = 32'd6
; 
32'd9522: dataIn1 = 32'd10
; 
32'd9523: dataIn1 = 32'd12
; 
32'd9524: dataIn1 = 32'd14
; 
32'd9525: dataIn1 = 32'd15
; 
32'd9526: dataIn1 = 32'd16
; 
32'd9527: dataIn1 = 32'd17
; 
32'd9528: dataIn1 = 32'd20
; 
32'd9529: dataIn1 = 32'd21
; 
32'd9530: dataIn1 = 32'd22
; 
32'd9531: dataIn1 = 32'd24
; 
32'd9532: dataIn1 = 32'd25
; 
32'd9533: dataIn1 = 32'd28
; 
32'd9534: dataIn1 = 32'd29
; 
32'd9535: dataIn1 = 32'd30
; 
32'd9536: dataIn1 = 32'd0
; 
32'd9537: dataIn1 = 32'd1
; 
32'd9538: dataIn1 = 32'd2
; 
32'd9539: dataIn1 = 32'd4
; 
32'd9540: dataIn1 = 32'd5
; 
32'd9541: dataIn1 = 32'd6
; 
32'd9542: dataIn1 = 32'd7
; 
32'd9543: dataIn1 = 32'd8
; 
32'd9544: dataIn1 = 32'd9
; 
32'd9545: dataIn1 = 32'd10
; 
32'd9546: dataIn1 = 32'd12
; 
32'd9547: dataIn1 = 32'd13
; 
32'd9548: dataIn1 = 32'd16
; 
32'd9549: dataIn1 = 32'd17
; 
32'd9550: dataIn1 = 32'd18
; 
32'd9551: dataIn1 = 32'd19
; 
32'd9552: dataIn1 = 32'd20
; 
32'd9553: dataIn1 = 32'd21
; 
32'd9554: dataIn1 = 32'd24
; 
32'd9555: dataIn1 = 32'd25
; 
32'd9556: dataIn1 = 32'd27
; 
32'd9557: dataIn1 = 32'd28
; 
32'd9558: dataIn1 = 32'd29
; 
32'd9559: dataIn1 = 32'd30
; 
32'd9560: dataIn1 = 32'd31
; 
32'd9561: dataIn1 = 32'd0
; 
32'd9562: dataIn1 = 32'd1
; 
32'd9563: dataIn1 = 32'd2
; 
32'd9564: dataIn1 = 32'd3
; 
32'd9565: dataIn1 = 32'd4
; 
32'd9566: dataIn1 = 32'd5
; 
32'd9567: dataIn1 = 32'd6
; 
32'd9568: dataIn1 = 32'd7
; 
32'd9569: dataIn1 = 32'd8
; 
32'd9570: dataIn1 = 32'd9
; 
32'd9571: dataIn1 = 32'd11
; 
32'd9572: dataIn1 = 32'd13
; 
32'd9573: dataIn1 = 32'd14
; 
32'd9574: dataIn1 = 32'd16
; 
32'd9575: dataIn1 = 32'd18
; 
32'd9576: dataIn1 = 32'd19
; 
32'd9577: dataIn1 = 32'd20
; 
32'd9578: dataIn1 = 32'd22
; 
32'd9579: dataIn1 = 32'd24
; 
32'd9580: dataIn1 = 32'd27
; 
32'd9581: dataIn1 = 32'd29
; 
32'd9582: dataIn1 = 32'd31
; 
32'd9583: dataIn1 = 32'd0
; 
32'd9584: dataIn1 = 32'd4
; 
32'd9585: dataIn1 = 32'd6
; 
32'd9586: dataIn1 = 32'd7
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd54; 
32'd3: dataIn2 = 32'd87; 
32'd4: dataIn2 = 32'd2; 
32'd5: dataIn2 = 32'd52; 
32'd6: dataIn2 = 32'd58; 
32'd7: dataIn2 = 32'd30; 
32'd8: dataIn2 = 32'd32; 
32'd9: dataIn2 = 32'd18; 
32'd10: dataIn2 = 32'd44; 
32'd11: dataIn2 = 32'd20; 
32'd12: dataIn2 = 32'd75; 
32'd13: dataIn2 = 32'd57; 
32'd14: dataIn2 = 32'd7; 
32'd15: dataIn2 = 32'd90; 
32'd16: dataIn2 = 32'd24; 
32'd17: dataIn2 = 32'd42; 
32'd18: dataIn2 = 32'd25; 
32'd19: dataIn2 = 32'd76; 
32'd20: dataIn2 = 32'd51; 
32'd21: dataIn2 = 32'd24; 
32'd22: dataIn2 = 32'd71; 
32'd23: dataIn2 = 32'd43; 
32'd24: dataIn2 = 32'd20; 
32'd25: dataIn2 = 32'd17; 
32'd26: dataIn2 = 32'd83; 
32'd27: dataIn2 = 32'd65; 
32'd28: dataIn2 = 32'd40; 
32'd29: dataIn2 = 32'd54; 
32'd30: dataIn2 = 32'd47; 
32'd31: dataIn2 = 32'd64; 
32'd32: dataIn2 = 32'd19; 
32'd33: dataIn2 = 32'd24; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd170: dataIn2 = 32'd78; 
32'd171: dataIn2 = 32'd52; 
32'd172: dataIn2 = 32'd69; 
32'd173: dataIn2 = 32'd1; 
32'd174: dataIn2 = 32'd69; 
32'd175: dataIn2 = 32'd7; 
32'd176: dataIn2 = 32'd87; 
32'd177: dataIn2 = 32'd14; 
32'd178: dataIn2 = 32'd68; 
32'd179: dataIn2 = 32'd48; 
32'd180: dataIn2 = 32'd34; 
32'd181: dataIn2 = 32'd82; 
32'd182: dataIn2 = 32'd56; 
32'd183: dataIn2 = 32'd58; 
32'd184: dataIn2 = 32'd38; 
32'd185: dataIn2 = 32'd88; 
32'd186: dataIn2 = 32'd77; 
32'd187: dataIn2 = 32'd51; 
32'd188: dataIn2 = 32'd21; 
32'd189: dataIn2 = 32'd47; 
32'd190: dataIn2 = 32'd74; 
32'd191: dataIn2 = 32'd70; 
32'd192: dataIn2 = 32'd55; 
32'd193: dataIn2 = 32'd44; 
32'd194: dataIn2 = 32'd70; 
32'd195: dataIn2 = 32'd68; 
32'd196: dataIn2 = 32'd45; 
32'd197: dataIn2 = 32'd20; 
32'd198: dataIn2 = 32'd85; 
32'd199: dataIn2 = 32'd23; 
32'd200: dataIn2 = 32'd45; 
32'd201: dataIn2 = 32'd70; 
32'd202: dataIn2 = 32'd89; 
32'd203: dataIn2 = 32'd45; 
32'd204: dataIn2 = 32'd45; 
32'd205: dataIn2 = 32'd67; 
32'd206: dataIn2 = 32'd98; 
32'd207: dataIn2 = 32'd46; 
32'd208: dataIn2 = 32'd31; 
32'd209: dataIn2 = 32'd51; 
32'd210: dataIn2 = 32'd0; 
32'd211: dataIn2 = 32'd91; 
32'd212: dataIn2 = 32'd59; 
32'd213: dataIn2 = 32'd78; 
32'd214: dataIn2 = 32'd8; 
32'd215: dataIn2 = 32'd82; 
32'd216: dataIn2 = 32'd96; 
32'd217: dataIn2 = 32'd74; 
32'd218: dataIn2 = 32'd94; 
32'd219: dataIn2 = 32'd38; 
32'd220: dataIn2 = 32'd61; 
32'd221: dataIn2 = 32'd93; 
32'd222: dataIn2 = 32'd33; 
32'd223: dataIn2 = 32'd96; 
32'd224: dataIn2 = 32'd32; 
32'd225: dataIn2 = 32'd2; 
32'd226: dataIn2 = 32'd66; 
32'd227: dataIn2 = 32'd69; 
32'd228: dataIn2 = 32'd29; 
32'd229: dataIn2 = 32'd9; 
32'd230: dataIn2 = 32'd72; 
32'd231: dataIn2 = 32'd100; 
32'd232: dataIn2 = 32'd64; 
32'd233: dataIn2 = 32'd4; 
32'd234: dataIn2 = 32'd58; 
32'd235: dataIn2 = 32'd23; 
32'd236: dataIn2 = 32'd83; 
32'd237: dataIn2 = 32'd45; 
32'd238: dataIn2 = 32'd70; 
32'd239: dataIn2 = 32'd84; 
32'd240: dataIn2 = 32'd26; 
32'd241: dataIn2 = 32'd74; 
32'd242: dataIn2 = 32'd52; 
32'd243: dataIn2 = 32'd26; 
32'd244: dataIn2 = 32'd69; 
32'd245: dataIn2 = 32'd29; 
32'd246: dataIn2 = 32'd76; 
32'd247: dataIn2 = 32'd69; 
32'd248: dataIn2 = 32'd56; 
32'd249: dataIn2 = 32'd70; 
32'd250: dataIn2 = 32'd36; 
32'd251: dataIn2 = 32'd47; 
32'd252: dataIn2 = 32'd76; 
32'd253: dataIn2 = 32'd51; 
32'd254: dataIn2 = 32'd30; 
32'd255: dataIn2 = 32'd91; 
32'd256: dataIn2 = 32'd58; 
32'd257: dataIn2 = 32'd59; 
32'd258: dataIn2 = 32'd53; 
32'd259: dataIn2 = 32'd74; 
32'd260: dataIn2 = 32'd52; 
32'd261: dataIn2 = 32'd89; 
32'd262: dataIn2 = 32'd51; 
32'd263: dataIn2 = 32'd27; 
32'd264: dataIn2 = 32'd57; 
32'd265: dataIn2 = 32'd39; 
32'd266: dataIn2 = 32'd69; 
32'd267: dataIn2 = 32'd0; 
32'd268: dataIn2 = 32'd16; 
32'd269: dataIn2 = 32'd98; 
32'd270: dataIn2 = 32'd42; 
32'd271: dataIn2 = 32'd32; 
32'd272: dataIn2 = 32'd51; 
32'd273: dataIn2 = 32'd62; 
32'd274: dataIn2 = 32'd57; 
32'd275: dataIn2 = 32'd65; 
32'd276: dataIn2 = 32'd16; 
32'd277: dataIn2 = 32'd67; 
32'd278: dataIn2 = 32'd0; 
32'd279: dataIn2 = 32'd83; 
32'd280: dataIn2 = 32'd97; 
32'd281: dataIn2 = 32'd55; 
32'd282: dataIn2 = 32'd63; 
32'd283: dataIn2 = 32'd14; 
32'd284: dataIn2 = 32'd25; 
32'd285: dataIn2 = 32'd32; 
32'd286: dataIn2 = 32'd85; 
32'd287: dataIn2 = 32'd18; 
32'd288: dataIn2 = 32'd95; 
32'd289: dataIn2 = 32'd6; 
32'd290: dataIn2 = 32'd54; 
32'd291: dataIn2 = 32'd78; 
32'd292: dataIn2 = 32'd47; 
32'd293: dataIn2 = 32'd97; 
32'd294: dataIn2 = 32'd78; 
32'd295: dataIn2 = 32'd97; 
32'd296: dataIn2 = 32'd42; 
32'd297: dataIn2 = 32'd10; 
32'd298: dataIn2 = 32'd31; 
32'd299: dataIn2 = 32'd97; 
32'd300: dataIn2 = 32'd99; 
32'd301: dataIn2 = 32'd80; 
32'd302: dataIn2 = 32'd28; 
32'd303: dataIn2 = 32'd26; 
32'd304: dataIn2 = 32'd20; 
32'd305: dataIn2 = 32'd66; 
32'd306: dataIn2 = 32'd28; 
32'd307: dataIn2 = 32'd53; 
32'd308: dataIn2 = 32'd74; 
32'd309: dataIn2 = 32'd52; 
32'd310: dataIn2 = 32'd91; 
32'd311: dataIn2 = 32'd23; 
32'd312: dataIn2 = 32'd69; 
32'd313: dataIn2 = 32'd60; 
32'd314: dataIn2 = 32'd71; 
32'd315: dataIn2 = 32'd73; 
32'd316: dataIn2 = 32'd8; 
32'd317: dataIn2 = 32'd55; 
32'd318: dataIn2 = 32'd2; 
32'd319: dataIn2 = 32'd9; 
32'd320: dataIn2 = 32'd87; 
32'd321: dataIn2 = 32'd93; 
32'd322: dataIn2 = 32'd45; 
32'd323: dataIn2 = 32'd68; 
32'd324: dataIn2 = 32'd62; 
32'd325: dataIn2 = 32'd63; 
32'd326: dataIn2 = 32'd17; 
32'd327: dataIn2 = 32'd31; 
32'd328: dataIn2 = 32'd79; 
32'd329: dataIn2 = 32'd57; 
32'd330: dataIn2 = 32'd34; 
32'd331: dataIn2 = 32'd91; 
32'd332: dataIn2 = 32'd0; 
32'd333: dataIn2 = 32'd29; 
32'd334: dataIn2 = 32'd25; 
32'd335: dataIn2 = 32'd63; 
32'd336: dataIn2 = 32'd85; 
32'd337: dataIn2 = 32'd9; 
32'd338: dataIn2 = 32'd25; 
32'd339: dataIn2 = 32'd19; 
32'd340: dataIn2 = 32'd65; 
32'd341: dataIn2 = 32'd56; 
32'd342: dataIn2 = 32'd54; 
32'd343: dataIn2 = 32'd67; 
32'd344: dataIn2 = 32'd93; 
32'd345: dataIn2 = 32'd92; 
32'd346: dataIn2 = 32'd94; 
32'd347: dataIn2 = 32'd90; 
32'd348: dataIn2 = 32'd15; 
32'd349: dataIn2 = 32'd56; 
32'd350: dataIn2 = 32'd25; 
32'd351: dataIn2 = 32'd58; 
32'd352: dataIn2 = 32'd68; 
32'd353: dataIn2 = 32'd48; 
32'd354: dataIn2 = 32'd39; 
32'd355: dataIn2 = 32'd23; 
32'd356: dataIn2 = 32'd33; 
32'd357: dataIn2 = 32'd36; 
32'd358: dataIn2 = 32'd58; 
32'd359: dataIn2 = 32'd35; 
32'd360: dataIn2 = 32'd72; 
32'd361: dataIn2 = 32'd35; 
32'd362: dataIn2 = 32'd75; 
32'd363: dataIn2 = 32'd66; 
32'd364: dataIn2 = 32'd53; 
32'd365: dataIn2 = 32'd91; 
32'd366: dataIn2 = 32'd77; 
32'd367: dataIn2 = 32'd26; 
32'd368: dataIn2 = 32'd71; 
32'd369: dataIn2 = 32'd95; 
32'd370: dataIn2 = 32'd78; 
32'd371: dataIn2 = 32'd87; 
32'd372: dataIn2 = 32'd42; 
32'd373: dataIn2 = 32'd76; 
32'd374: dataIn2 = 32'd100; 
32'd375: dataIn2 = 32'd84; 
32'd376: dataIn2 = 32'd49; 
32'd377: dataIn2 = 32'd79; 
32'd378: dataIn2 = 32'd62; 
32'd379: dataIn2 = 32'd32; 
32'd380: dataIn2 = 32'd1; 
32'd381: dataIn2 = 32'd81; 
32'd382: dataIn2 = 32'd28; 
32'd383: dataIn2 = 32'd17; 
32'd384: dataIn2 = 32'd77; 
32'd385: dataIn2 = 32'd75; 
32'd386: dataIn2 = 32'd11; 
32'd387: dataIn2 = 32'd76; 
32'd388: dataIn2 = 32'd58; 
32'd389: dataIn2 = 32'd8; 
32'd390: dataIn2 = 32'd61; 
32'd391: dataIn2 = 32'd50; 
32'd392: dataIn2 = 32'd68; 
32'd393: dataIn2 = 32'd55; 
32'd394: dataIn2 = 32'd15; 
32'd395: dataIn2 = 32'd68; 
32'd396: dataIn2 = 32'd99; 
32'd397: dataIn2 = 32'd35; 
32'd398: dataIn2 = 32'd59; 
32'd399: dataIn2 = 32'd26; 
32'd400: dataIn2 = 32'd65; 
32'd401: dataIn2 = 32'd82; 
32'd402: dataIn2 = 32'd15; 
32'd403: dataIn2 = 32'd59; 
32'd404: dataIn2 = 32'd19; 
32'd405: dataIn2 = 32'd74; 
32'd406: dataIn2 = 32'd39; 
32'd407: dataIn2 = 32'd52; 
32'd408: dataIn2 = 32'd1; 
32'd409: dataIn2 = 32'd50; 
32'd410: dataIn2 = 32'd22; 
32'd411: dataIn2 = 32'd80; 
32'd412: dataIn2 = 32'd86; 
32'd413: dataIn2 = 32'd26; 
32'd414: dataIn2 = 32'd22; 
32'd415: dataIn2 = 32'd68; 
32'd416: dataIn2 = 32'd20; 
32'd417: dataIn2 = 32'd10; 
32'd418: dataIn2 = 32'd50; 
32'd419: dataIn2 = 32'd12; 
32'd420: dataIn2 = 32'd85; 
32'd421: dataIn2 = 32'd84; 
32'd422: dataIn2 = 32'd1; 
32'd423: dataIn2 = 32'd16; 
32'd424: dataIn2 = 32'd48; 
32'd425: dataIn2 = 32'd38; 
32'd426: dataIn2 = 32'd33; 
32'd427: dataIn2 = 32'd46; 
32'd428: dataIn2 = 32'd4; 
32'd429: dataIn2 = 32'd79; 
32'd430: dataIn2 = 32'd66; 
32'd431: dataIn2 = 32'd65; 
32'd432: dataIn2 = 32'd50; 
32'd433: dataIn2 = 32'd89; 
32'd434: dataIn2 = 32'd22; 
32'd435: dataIn2 = 32'd83; 
32'd436: dataIn2 = 32'd14; 
32'd437: dataIn2 = 32'd59; 
32'd438: dataIn2 = 32'd46; 
32'd439: dataIn2 = 32'd54; 
32'd440: dataIn2 = 32'd84; 
32'd441: dataIn2 = 32'd88; 
32'd442: dataIn2 = 32'd99; 
32'd443: dataIn2 = 32'd32; 
32'd444: dataIn2 = 32'd9; 
32'd445: dataIn2 = 32'd96; 
32'd446: dataIn2 = 32'd33; 
32'd447: dataIn2 = 32'd83; 
32'd448: dataIn2 = 32'd47; 
32'd449: dataIn2 = 32'd88; 
32'd450: dataIn2 = 32'd20; 
32'd451: dataIn2 = 32'd60; 
32'd452: dataIn2 = 32'd6; 
32'd453: dataIn2 = 32'd1; 
32'd454: dataIn2 = 32'd46; 
32'd455: dataIn2 = 32'd13; 
32'd456: dataIn2 = 32'd84; 
32'd457: dataIn2 = 32'd41; 
32'd458: dataIn2 = 32'd85; 
32'd459: dataIn2 = 32'd81; 
32'd460: dataIn2 = 32'd82; 
32'd461: dataIn2 = 32'd89; 
32'd462: dataIn2 = 32'd49; 
32'd463: dataIn2 = 32'd62; 
32'd464: dataIn2 = 32'd78; 
32'd465: dataIn2 = 32'd1; 
32'd466: dataIn2 = 32'd28; 
32'd467: dataIn2 = 32'd98; 
32'd468: dataIn2 = 32'd65; 
32'd469: dataIn2 = 32'd100; 
32'd470: dataIn2 = 32'd69; 
32'd471: dataIn2 = 32'd66; 
32'd472: dataIn2 = 32'd31; 
32'd473: dataIn2 = 32'd60; 
32'd474: dataIn2 = 32'd36; 
32'd475: dataIn2 = 32'd3; 
32'd476: dataIn2 = 32'd29; 
32'd477: dataIn2 = 32'd17; 
32'd478: dataIn2 = 32'd4; 
32'd479: dataIn2 = 32'd75; 
32'd480: dataIn2 = 32'd2; 
32'd481: dataIn2 = 32'd48; 
32'd482: dataIn2 = 32'd41; 
32'd483: dataIn2 = 32'd29; 
32'd484: dataIn2 = 32'd43; 
32'd485: dataIn2 = 32'd83; 
32'd486: dataIn2 = 32'd67; 
32'd487: dataIn2 = 32'd56; 
32'd488: dataIn2 = 32'd0; 
32'd489: dataIn2 = 32'd27; 
32'd490: dataIn2 = 32'd94; 
32'd491: dataIn2 = 32'd19; 
32'd492: dataIn2 = 32'd28; 
32'd493: dataIn2 = 32'd80; 
32'd494: dataIn2 = 32'd72; 
32'd495: dataIn2 = 32'd9; 
32'd496: dataIn2 = 32'd92; 
32'd497: dataIn2 = 32'd72; 
32'd498: dataIn2 = 32'd44; 
32'd499: dataIn2 = 32'd18; 
32'd500: dataIn2 = 32'd84; 
32'd501: dataIn2 = 32'd77; 
32'd502: dataIn2 = 32'd100; 
32'd503: dataIn2 = 32'd22; 
32'd504: dataIn2 = 32'd94; 
32'd505: dataIn2 = 32'd12; 
32'd506: dataIn2 = 32'd62; 
32'd507: dataIn2 = 32'd85; 
32'd508: dataIn2 = 32'd86; 
32'd509: dataIn2 = 32'd80; 
32'd510: dataIn2 = 32'd85; 
32'd511: dataIn2 = 32'd64; 
32'd512: dataIn2 = 32'd16; 
32'd513: dataIn2 = 32'd68; 
32'd514: dataIn2 = 32'd33; 
32'd515: dataIn2 = 32'd99; 
32'd516: dataIn2 = 32'd38; 
32'd517: dataIn2 = 32'd91; 
32'd518: dataIn2 = 32'd29; 
32'd519: dataIn2 = 32'd50; 
32'd520: dataIn2 = 32'd35; 
32'd521: dataIn2 = 32'd41; 
32'd522: dataIn2 = 32'd4; 
32'd523: dataIn2 = 32'd0; 
32'd524: dataIn2 = 32'd7; 
32'd525: dataIn2 = 32'd17; 
32'd526: dataIn2 = 32'd88; 
32'd527: dataIn2 = 32'd39; 
32'd528: dataIn2 = 32'd28; 
32'd529: dataIn2 = 32'd67; 
32'd530: dataIn2 = 32'd77; 
32'd531: dataIn2 = 32'd86; 
32'd532: dataIn2 = 32'd96; 
32'd533: dataIn2 = 32'd20; 
32'd534: dataIn2 = 32'd68; 
32'd535: dataIn2 = 32'd8; 
32'd536: dataIn2 = 32'd80; 
32'd537: dataIn2 = 32'd62; 
32'd538: dataIn2 = 32'd46; 
32'd539: dataIn2 = 32'd11; 
32'd540: dataIn2 = 32'd12; 
32'd541: dataIn2 = 32'd87; 
32'd542: dataIn2 = 32'd5; 
32'd543: dataIn2 = 32'd71; 
32'd544: dataIn2 = 32'd0; 
32'd545: dataIn2 = 32'd41; 
32'd546: dataIn2 = 32'd3; 
32'd547: dataIn2 = 32'd73; 
32'd548: dataIn2 = 32'd50; 
32'd549: dataIn2 = 32'd36; 
32'd550: dataIn2 = 32'd52; 
32'd551: dataIn2 = 32'd40; 
32'd552: dataIn2 = 32'd92; 
32'd553: dataIn2 = 32'd90; 
32'd554: dataIn2 = 32'd3; 
32'd555: dataIn2 = 32'd99; 
32'd556: dataIn2 = 32'd56; 
32'd557: dataIn2 = 32'd68; 
32'd558: dataIn2 = 32'd92; 
32'd559: dataIn2 = 32'd52; 
32'd560: dataIn2 = 32'd87; 
32'd561: dataIn2 = 32'd27; 
32'd562: dataIn2 = 32'd52; 
32'd563: dataIn2 = 32'd59; 
32'd564: dataIn2 = 32'd14; 
32'd565: dataIn2 = 32'd5; 
32'd566: dataIn2 = 32'd37; 
32'd567: dataIn2 = 32'd39; 
32'd568: dataIn2 = 32'd33; 
32'd569: dataIn2 = 32'd79; 
32'd570: dataIn2 = 32'd88; 
32'd571: dataIn2 = 32'd37; 
32'd572: dataIn2 = 32'd7; 
32'd573: dataIn2 = 32'd15; 
32'd574: dataIn2 = 32'd62; 
32'd575: dataIn2 = 32'd5; 
32'd576: dataIn2 = 32'd95; 
32'd577: dataIn2 = 32'd57; 
32'd578: dataIn2 = 32'd3; 
32'd579: dataIn2 = 32'd96; 
32'd580: dataIn2 = 32'd92; 
32'd581: dataIn2 = 32'd31; 
32'd582: dataIn2 = 32'd52; 
32'd583: dataIn2 = 32'd35; 
32'd584: dataIn2 = 32'd88; 
32'd585: dataIn2 = 32'd80; 
32'd586: dataIn2 = 32'd89; 
32'd587: dataIn2 = 32'd45; 
32'd588: dataIn2 = 32'd44; 
32'd589: dataIn2 = 32'd83; 
32'd590: dataIn2 = 32'd61; 
32'd591: dataIn2 = 32'd73; 
32'd592: dataIn2 = 32'd9; 
32'd593: dataIn2 = 32'd22; 
32'd594: dataIn2 = 32'd42; 
32'd595: dataIn2 = 32'd22; 
32'd596: dataIn2 = 32'd8; 
32'd597: dataIn2 = 32'd78; 
32'd598: dataIn2 = 32'd4; 
32'd599: dataIn2 = 32'd51; 
32'd600: dataIn2 = 32'd10; 
32'd601: dataIn2 = 32'd48; 
32'd602: dataIn2 = 32'd12; 
32'd603: dataIn2 = 32'd94; 
32'd604: dataIn2 = 32'd44; 
32'd605: dataIn2 = 32'd23; 
32'd606: dataIn2 = 32'd19; 
32'd607: dataIn2 = 32'd46; 
32'd608: dataIn2 = 32'd80; 
32'd609: dataIn2 = 32'd73; 
32'd610: dataIn2 = 32'd56; 
32'd611: dataIn2 = 32'd92; 
32'd612: dataIn2 = 32'd69; 
32'd613: dataIn2 = 32'd71; 
32'd614: dataIn2 = 32'd22; 
32'd615: dataIn2 = 32'd42; 
32'd616: dataIn2 = 32'd62; 
32'd617: dataIn2 = 32'd41; 
32'd618: dataIn2 = 32'd33; 
32'd619: dataIn2 = 32'd95; 
32'd620: dataIn2 = 32'd15; 
32'd621: dataIn2 = 32'd42; 
32'd622: dataIn2 = 32'd79; 
32'd623: dataIn2 = 32'd66; 
32'd624: dataIn2 = 32'd60; 
32'd625: dataIn2 = 32'd11; 
32'd626: dataIn2 = 32'd5; 
32'd627: dataIn2 = 32'd88; 
32'd628: dataIn2 = 32'd92; 
32'd629: dataIn2 = 32'd95; 
32'd630: dataIn2 = 32'd46; 
32'd631: dataIn2 = 32'd49; 
32'd632: dataIn2 = 32'd68; 
32'd633: dataIn2 = 32'd23; 
32'd634: dataIn2 = 32'd57; 
32'd635: dataIn2 = 32'd71; 
32'd636: dataIn2 = 32'd97; 
32'd637: dataIn2 = 32'd66; 
32'd638: dataIn2 = 32'd6; 
32'd639: dataIn2 = 32'd5; 
32'd640: dataIn2 = 32'd74; 
32'd641: dataIn2 = 32'd74; 
32'd642: dataIn2 = 32'd44; 
32'd643: dataIn2 = 32'd38; 
32'd644: dataIn2 = 32'd24; 
32'd645: dataIn2 = 32'd92; 
32'd646: dataIn2 = 32'd80; 
32'd647: dataIn2 = 32'd42; 
32'd648: dataIn2 = 32'd0; 
32'd649: dataIn2 = 32'd32; 
32'd650: dataIn2 = 32'd31; 
32'd651: dataIn2 = 32'd78; 
32'd652: dataIn2 = 32'd81; 
32'd653: dataIn2 = 32'd50; 
32'd654: dataIn2 = 32'd7; 
32'd655: dataIn2 = 32'd17; 
32'd656: dataIn2 = 32'd16; 
32'd657: dataIn2 = 32'd92; 
32'd658: dataIn2 = 32'd95; 
32'd659: dataIn2 = 32'd50; 
32'd660: dataIn2 = 32'd9; 
32'd661: dataIn2 = 32'd87; 
32'd662: dataIn2 = 32'd88; 
32'd663: dataIn2 = 32'd32; 
32'd664: dataIn2 = 32'd28; 
32'd665: dataIn2 = 32'd34; 
32'd666: dataIn2 = 32'd16; 
32'd667: dataIn2 = 32'd25; 
32'd668: dataIn2 = 32'd80; 
32'd669: dataIn2 = 32'd24; 
32'd670: dataIn2 = 32'd42; 
32'd671: dataIn2 = 32'd22; 
32'd672: dataIn2 = 32'd81; 
32'd673: dataIn2 = 32'd22; 
32'd674: dataIn2 = 32'd17; 
32'd675: dataIn2 = 32'd75; 
32'd676: dataIn2 = 32'd3; 
32'd677: dataIn2 = 32'd6; 
32'd678: dataIn2 = 32'd50; 
32'd679: dataIn2 = 32'd10; 
32'd680: dataIn2 = 32'd52; 
32'd681: dataIn2 = 32'd80; 
32'd682: dataIn2 = 32'd53; 
32'd683: dataIn2 = 32'd30; 
32'd684: dataIn2 = 32'd29; 
32'd685: dataIn2 = 32'd96; 
32'd686: dataIn2 = 32'd11; 
32'd687: dataIn2 = 32'd62; 
32'd688: dataIn2 = 32'd91; 
32'd689: dataIn2 = 32'd30; 
32'd690: dataIn2 = 32'd21; 
32'd691: dataIn2 = 32'd85; 
32'd692: dataIn2 = 32'd49; 
32'd693: dataIn2 = 32'd55; 
32'd694: dataIn2 = 32'd48; 
32'd695: dataIn2 = 32'd34; 
32'd696: dataIn2 = 32'd78; 
32'd697: dataIn2 = 32'd67; 
32'd698: dataIn2 = 32'd33; 
32'd699: dataIn2 = 32'd11; 
32'd700: dataIn2 = 32'd59; 
32'd701: dataIn2 = 32'd21; 
32'd702: dataIn2 = 32'd65; 
32'd703: dataIn2 = 32'd49; 
32'd704: dataIn2 = 32'd37; 
32'd705: dataIn2 = 32'd80; 
32'd706: dataIn2 = 32'd30; 
32'd707: dataIn2 = 32'd26; 
32'd708: dataIn2 = 32'd28; 
32'd709: dataIn2 = 32'd32; 
32'd710: dataIn2 = 32'd66; 
32'd711: dataIn2 = 32'd99; 
32'd712: dataIn2 = 32'd28; 
32'd713: dataIn2 = 32'd13; 
32'd714: dataIn2 = 32'd73; 
32'd715: dataIn2 = 32'd40; 
32'd716: dataIn2 = 32'd68; 
32'd717: dataIn2 = 32'd49; 
32'd718: dataIn2 = 32'd62; 
32'd719: dataIn2 = 32'd48; 
32'd720: dataIn2 = 32'd5; 
32'd721: dataIn2 = 32'd17; 
32'd722: dataIn2 = 32'd6; 
32'd723: dataIn2 = 32'd95; 
32'd724: dataIn2 = 32'd27; 
32'd725: dataIn2 = 32'd42; 
32'd726: dataIn2 = 32'd36; 
32'd727: dataIn2 = 32'd62; 
32'd728: dataIn2 = 32'd59; 
32'd729: dataIn2 = 32'd8; 
32'd730: dataIn2 = 32'd85; 
32'd731: dataIn2 = 32'd86; 
32'd732: dataIn2 = 32'd38; 
32'd733: dataIn2 = 32'd28; 
32'd734: dataIn2 = 32'd7; 
32'd735: dataIn2 = 32'd83; 
32'd736: dataIn2 = 32'd97; 
32'd737: dataIn2 = 32'd16; 
32'd738: dataIn2 = 32'd42; 
32'd739: dataIn2 = 32'd39; 
32'd740: dataIn2 = 32'd43; 
32'd741: dataIn2 = 32'd85; 
32'd742: dataIn2 = 32'd32; 
32'd743: dataIn2 = 32'd13; 
32'd744: dataIn2 = 32'd55; 
32'd745: dataIn2 = 32'd13; 
32'd746: dataIn2 = 32'd2; 
32'd747: dataIn2 = 32'd71; 
32'd748: dataIn2 = 32'd85; 
32'd749: dataIn2 = 32'd33; 
32'd750: dataIn2 = 32'd55; 
32'd751: dataIn2 = 32'd32; 
32'd752: dataIn2 = 32'd9; 
32'd753: dataIn2 = 32'd62; 
32'd754: dataIn2 = 32'd12; 
32'd755: dataIn2 = 32'd2; 
32'd756: dataIn2 = 32'd98; 
32'd757: dataIn2 = 32'd42; 
32'd758: dataIn2 = 32'd69; 
32'd759: dataIn2 = 32'd95; 
32'd760: dataIn2 = 32'd30; 
32'd761: dataIn2 = 32'd92; 
32'd762: dataIn2 = 32'd29; 
32'd763: dataIn2 = 32'd50; 
32'd764: dataIn2 = 32'd42; 
32'd765: dataIn2 = 32'd58; 
32'd766: dataIn2 = 32'd20; 
32'd767: dataIn2 = 32'd66; 
32'd768: dataIn2 = 32'd9; 
32'd769: dataIn2 = 32'd64; 
32'd770: dataIn2 = 32'd35; 
32'd771: dataIn2 = 32'd83; 
32'd772: dataIn2 = 32'd20; 
32'd773: dataIn2 = 32'd61; 
32'd774: dataIn2 = 32'd53; 
32'd775: dataIn2 = 32'd91; 
32'd776: dataIn2 = 32'd93; 
32'd777: dataIn2 = 32'd59; 
32'd778: dataIn2 = 32'd91; 
32'd779: dataIn2 = 32'd65; 
32'd780: dataIn2 = 32'd53; 
32'd781: dataIn2 = 32'd52; 
32'd782: dataIn2 = 32'd3; 
32'd783: dataIn2 = 32'd29; 
32'd784: dataIn2 = 32'd90; 
32'd785: dataIn2 = 32'd11; 
32'd786: dataIn2 = 32'd74; 
32'd787: dataIn2 = 32'd48; 
32'd788: dataIn2 = 32'd83; 
32'd789: dataIn2 = 32'd91; 
32'd790: dataIn2 = 32'd32; 
32'd791: dataIn2 = 32'd44; 
32'd792: dataIn2 = 32'd32; 
32'd793: dataIn2 = 32'd85; 
32'd794: dataIn2 = 32'd25; 
32'd795: dataIn2 = 32'd75; 
32'd796: dataIn2 = 32'd72; 
32'd797: dataIn2 = 32'd19; 
32'd798: dataIn2 = 32'd54; 
32'd799: dataIn2 = 32'd21; 
32'd800: dataIn2 = 32'd33; 
32'd801: dataIn2 = 32'd21; 
32'd802: dataIn2 = 32'd25; 
32'd803: dataIn2 = 32'd57; 
32'd804: dataIn2 = 32'd5; 
32'd805: dataIn2 = 32'd14; 
32'd806: dataIn2 = 32'd58; 
32'd807: dataIn2 = 32'd40; 
32'd808: dataIn2 = 32'd68; 
32'd809: dataIn2 = 32'd80; 
32'd810: dataIn2 = 32'd1; 
32'd811: dataIn2 = 32'd96; 
32'd812: dataIn2 = 32'd20; 
32'd813: dataIn2 = 32'd52; 
32'd814: dataIn2 = 32'd32; 
32'd815: dataIn2 = 32'd78; 
32'd816: dataIn2 = 32'd21; 
32'd817: dataIn2 = 32'd77; 
32'd818: dataIn2 = 32'd47; 
32'd819: dataIn2 = 32'd47; 
32'd820: dataIn2 = 32'd49; 
32'd821: dataIn2 = 32'd30; 
32'd822: dataIn2 = 32'd24; 
32'd823: dataIn2 = 32'd43; 
32'd824: dataIn2 = 32'd84; 
32'd825: dataIn2 = 32'd41; 
32'd826: dataIn2 = 32'd16; 
32'd827: dataIn2 = 32'd70; 
32'd828: dataIn2 = 32'd100; 
32'd829: dataIn2 = 32'd19; 
32'd830: dataIn2 = 32'd11; 
32'd831: dataIn2 = 32'd95; 
32'd832: dataIn2 = 32'd78; 
32'd833: dataIn2 = 32'd65; 
32'd834: dataIn2 = 32'd61; 
32'd835: dataIn2 = 32'd94; 
32'd836: dataIn2 = 32'd59; 
32'd837: dataIn2 = 32'd37; 
32'd838: dataIn2 = 32'd57; 
32'd839: dataIn2 = 32'd18; 
32'd840: dataIn2 = 32'd63; 
32'd841: dataIn2 = 32'd57; 
32'd842: dataIn2 = 32'd35; 
32'd843: dataIn2 = 32'd10; 
32'd844: dataIn2 = 32'd56; 
32'd845: dataIn2 = 32'd93; 
32'd846: dataIn2 = 32'd70; 
32'd847: dataIn2 = 32'd19; 
32'd848: dataIn2 = 32'd20; 
32'd849: dataIn2 = 32'd53; 
32'd850: dataIn2 = 32'd83; 
32'd851: dataIn2 = 32'd49; 
32'd852: dataIn2 = 32'd25; 
32'd853: dataIn2 = 32'd15; 
32'd854: dataIn2 = 32'd76; 
32'd855: dataIn2 = 32'd24; 
32'd856: dataIn2 = 32'd15; 
32'd857: dataIn2 = 32'd76; 
32'd858: dataIn2 = 32'd73; 
32'd859: dataIn2 = 32'd94; 
32'd860: dataIn2 = 32'd31; 
32'd861: dataIn2 = 32'd76; 
32'd862: dataIn2 = 32'd13; 
32'd863: dataIn2 = 32'd64; 
32'd864: dataIn2 = 32'd60; 
32'd865: dataIn2 = 32'd19; 
32'd866: dataIn2 = 32'd31; 
32'd867: dataIn2 = 32'd7; 
32'd868: dataIn2 = 32'd23; 
32'd869: dataIn2 = 32'd24; 
32'd870: dataIn2 = 32'd41; 
32'd871: dataIn2 = 32'd46; 
32'd872: dataIn2 = 32'd70; 
32'd873: dataIn2 = 32'd29; 
32'd874: dataIn2 = 32'd2; 
32'd875: dataIn2 = 32'd3; 
32'd876: dataIn2 = 32'd96; 
32'd877: dataIn2 = 32'd36; 
32'd878: dataIn2 = 32'd72; 
32'd879: dataIn2 = 32'd66; 
32'd880: dataIn2 = 32'd95; 
32'd881: dataIn2 = 32'd40; 
32'd882: dataIn2 = 32'd20; 
32'd883: dataIn2 = 32'd17; 
32'd884: dataIn2 = 32'd43; 
32'd885: dataIn2 = 32'd28; 
32'd886: dataIn2 = 32'd44; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_32_30.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
