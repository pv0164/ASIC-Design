//32x32 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 614 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd170 ; 
  wdata_col_base = 32'd7840 ; 
  row_base = 32'd84540 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #12460; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd84540: dataIn1 = 32'd0
; 
32'd84541: dataIn1 = 32'd14
; 
32'd84542: dataIn1 = 32'd29
; 
32'd84543: dataIn1 = 32'd47
; 
32'd84544: dataIn1 = 32'd63
; 
32'd84545: dataIn1 = 32'd82
; 
32'd84546: dataIn1 = 32'd99
; 
32'd84547: dataIn1 = 32'd116
; 
32'd84548: dataIn1 = 32'd132
; 
32'd84549: dataIn1 = 32'd146
; 
32'd84550: dataIn1 = 32'd166
; 
32'd84551: dataIn1 = 32'd185
; 
32'd84552: dataIn1 = 32'd206
; 
32'd84553: dataIn1 = 32'd231
; 
32'd84554: dataIn1 = 32'd248
; 
32'd84555: dataIn1 = 32'd270
; 
32'd84556: dataIn1 = 32'd291
; 
32'd84557: dataIn1 = 32'd309
; 
32'd84558: dataIn1 = 32'd330
; 
32'd84559: dataIn1 = 32'd351
; 
32'd84560: dataIn1 = 32'd364
; 
32'd84561: dataIn1 = 32'd381
; 
32'd84562: dataIn1 = 32'd399
; 
32'd84563: dataIn1 = 32'd417
; 
32'd84564: dataIn1 = 32'd434
; 
32'd84565: dataIn1 = 32'd454
; 
32'd84566: dataIn1 = 32'd475
; 
32'd84567: dataIn1 = 32'd494
; 
32'd84568: dataIn1 = 32'd509
; 
32'd84569: dataIn1 = 32'd533
; 
32'd84570: dataIn1 = 32'd553
; 
32'd84571: dataIn1 = 32'd572
; 
32'd84572: dataIn1 = 32'd586
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd7840: dataIn1 = 32'd0
; 
32'd7841: dataIn1 = 32'd14
; 
32'd7842: dataIn1 = 32'd29
; 
32'd7843: dataIn1 = 32'd47
; 
32'd7844: dataIn1 = 32'd63
; 
32'd7845: dataIn1 = 32'd82
; 
32'd7846: dataIn1 = 32'd99
; 
32'd7847: dataIn1 = 32'd116
; 
32'd7848: dataIn1 = 32'd132
; 
32'd7849: dataIn1 = 32'd146
; 
32'd7850: dataIn1 = 32'd166
; 
32'd7851: dataIn1 = 32'd185
; 
32'd7852: dataIn1 = 32'd206
; 
32'd7853: dataIn1 = 32'd231
; 
32'd7854: dataIn1 = 32'd248
; 
32'd7855: dataIn1 = 32'd270
; 
32'd7856: dataIn1 = 32'd291
; 
32'd7857: dataIn1 = 32'd309
; 
32'd7858: dataIn1 = 32'd330
; 
32'd7859: dataIn1 = 32'd351
; 
32'd7860: dataIn1 = 32'd364
; 
32'd7861: dataIn1 = 32'd381
; 
32'd7862: dataIn1 = 32'd399
; 
32'd7863: dataIn1 = 32'd417
; 
32'd7864: dataIn1 = 32'd434
; 
32'd7865: dataIn1 = 32'd454
; 
32'd7866: dataIn1 = 32'd475
; 
32'd7867: dataIn1 = 32'd494
; 
32'd7868: dataIn1 = 32'd509
; 
32'd7869: dataIn1 = 32'd533
; 
32'd7870: dataIn1 = 32'd553
; 
32'd7871: dataIn1 = 32'd572
; 
32'd7872: dataIn1 = 32'd586
; 
32'd7873: dataIn1 = 32'd0
; 
32'd7874: dataIn1 = 32'd1
; 
32'd7875: dataIn1 = 32'd6
; 
32'd7876: dataIn1 = 32'd7
; 
32'd7877: dataIn1 = 32'd8
; 
32'd7878: dataIn1 = 32'd10
; 
32'd7879: dataIn1 = 32'd11
; 
32'd7880: dataIn1 = 32'd20
; 
32'd7881: dataIn1 = 32'd21
; 
32'd7882: dataIn1 = 32'd22
; 
32'd7883: dataIn1 = 32'd25
; 
32'd7884: dataIn1 = 32'd26
; 
32'd7885: dataIn1 = 32'd27
; 
32'd7886: dataIn1 = 32'd31
; 
32'd7887: dataIn1 = 32'd2
; 
32'd7888: dataIn1 = 32'd4
; 
32'd7889: dataIn1 = 32'd5
; 
32'd7890: dataIn1 = 32'd9
; 
32'd7891: dataIn1 = 32'd10
; 
32'd7892: dataIn1 = 32'd14
; 
32'd7893: dataIn1 = 32'd15
; 
32'd7894: dataIn1 = 32'd16
; 
32'd7895: dataIn1 = 32'd17
; 
32'd7896: dataIn1 = 32'd18
; 
32'd7897: dataIn1 = 32'd20
; 
32'd7898: dataIn1 = 32'd21
; 
32'd7899: dataIn1 = 32'd22
; 
32'd7900: dataIn1 = 32'd24
; 
32'd7901: dataIn1 = 32'd26
; 
32'd7902: dataIn1 = 32'd1
; 
32'd7903: dataIn1 = 32'd2
; 
32'd7904: dataIn1 = 32'd3
; 
32'd7905: dataIn1 = 32'd7
; 
32'd7906: dataIn1 = 32'd8
; 
32'd7907: dataIn1 = 32'd11
; 
32'd7908: dataIn1 = 32'd13
; 
32'd7909: dataIn1 = 32'd14
; 
32'd7910: dataIn1 = 32'd16
; 
32'd7911: dataIn1 = 32'd17
; 
32'd7912: dataIn1 = 32'd19
; 
32'd7913: dataIn1 = 32'd20
; 
32'd7914: dataIn1 = 32'd23
; 
32'd7915: dataIn1 = 32'd24
; 
32'd7916: dataIn1 = 32'd27
; 
32'd7917: dataIn1 = 32'd29
; 
32'd7918: dataIn1 = 32'd30
; 
32'd7919: dataIn1 = 32'd31
; 
32'd7920: dataIn1 = 32'd1
; 
32'd7921: dataIn1 = 32'd2
; 
32'd7922: dataIn1 = 32'd6
; 
32'd7923: dataIn1 = 32'd7
; 
32'd7924: dataIn1 = 32'd8
; 
32'd7925: dataIn1 = 32'd10
; 
32'd7926: dataIn1 = 32'd14
; 
32'd7927: dataIn1 = 32'd15
; 
32'd7928: dataIn1 = 32'd16
; 
32'd7929: dataIn1 = 32'd17
; 
32'd7930: dataIn1 = 32'd18
; 
32'd7931: dataIn1 = 32'd19
; 
32'd7932: dataIn1 = 32'd20
; 
32'd7933: dataIn1 = 32'd27
; 
32'd7934: dataIn1 = 32'd29
; 
32'd7935: dataIn1 = 32'd31
; 
32'd7936: dataIn1 = 32'd0
; 
32'd7937: dataIn1 = 32'd1
; 
32'd7938: dataIn1 = 32'd4
; 
32'd7939: dataIn1 = 32'd5
; 
32'd7940: dataIn1 = 32'd7
; 
32'd7941: dataIn1 = 32'd8
; 
32'd7942: dataIn1 = 32'd11
; 
32'd7943: dataIn1 = 32'd12
; 
32'd7944: dataIn1 = 32'd13
; 
32'd7945: dataIn1 = 32'd14
; 
32'd7946: dataIn1 = 32'd15
; 
32'd7947: dataIn1 = 32'd16
; 
32'd7948: dataIn1 = 32'd17
; 
32'd7949: dataIn1 = 32'd19
; 
32'd7950: dataIn1 = 32'd22
; 
32'd7951: dataIn1 = 32'd24
; 
32'd7952: dataIn1 = 32'd25
; 
32'd7953: dataIn1 = 32'd28
; 
32'd7954: dataIn1 = 32'd30
; 
32'd7955: dataIn1 = 32'd0
; 
32'd7956: dataIn1 = 32'd2
; 
32'd7957: dataIn1 = 32'd4
; 
32'd7958: dataIn1 = 32'd5
; 
32'd7959: dataIn1 = 32'd8
; 
32'd7960: dataIn1 = 32'd12
; 
32'd7961: dataIn1 = 32'd14
; 
32'd7962: dataIn1 = 32'd17
; 
32'd7963: dataIn1 = 32'd18
; 
32'd7964: dataIn1 = 32'd19
; 
32'd7965: dataIn1 = 32'd22
; 
32'd7966: dataIn1 = 32'd24
; 
32'd7967: dataIn1 = 32'd25
; 
32'd7968: dataIn1 = 32'd26
; 
32'd7969: dataIn1 = 32'd28
; 
32'd7970: dataIn1 = 32'd29
; 
32'd7971: dataIn1 = 32'd31
; 
32'd7972: dataIn1 = 32'd2
; 
32'd7973: dataIn1 = 32'd3
; 
32'd7974: dataIn1 = 32'd4
; 
32'd7975: dataIn1 = 32'd5
; 
32'd7976: dataIn1 = 32'd9
; 
32'd7977: dataIn1 = 32'd10
; 
32'd7978: dataIn1 = 32'd11
; 
32'd7979: dataIn1 = 32'd16
; 
32'd7980: dataIn1 = 32'd18
; 
32'd7981: dataIn1 = 32'd19
; 
32'd7982: dataIn1 = 32'd21
; 
32'd7983: dataIn1 = 32'd22
; 
32'd7984: dataIn1 = 32'd23
; 
32'd7985: dataIn1 = 32'd25
; 
32'd7986: dataIn1 = 32'd26
; 
32'd7987: dataIn1 = 32'd29
; 
32'd7988: dataIn1 = 32'd31
; 
32'd7989: dataIn1 = 32'd0
; 
32'd7990: dataIn1 = 32'd1
; 
32'd7991: dataIn1 = 32'd5
; 
32'd7992: dataIn1 = 32'd6
; 
32'd7993: dataIn1 = 32'd8
; 
32'd7994: dataIn1 = 32'd9
; 
32'd7995: dataIn1 = 32'd14
; 
32'd7996: dataIn1 = 32'd15
; 
32'd7997: dataIn1 = 32'd17
; 
32'd7998: dataIn1 = 32'd19
; 
32'd7999: dataIn1 = 32'd24
; 
32'd8000: dataIn1 = 32'd25
; 
32'd8001: dataIn1 = 32'd26
; 
32'd8002: dataIn1 = 32'd27
; 
32'd8003: dataIn1 = 32'd30
; 
32'd8004: dataIn1 = 32'd31
; 
32'd8005: dataIn1 = 32'd1
; 
32'd8006: dataIn1 = 32'd4
; 
32'd8007: dataIn1 = 32'd11
; 
32'd8008: dataIn1 = 32'd12
; 
32'd8009: dataIn1 = 32'd13
; 
32'd8010: dataIn1 = 32'd14
; 
32'd8011: dataIn1 = 32'd15
; 
32'd8012: dataIn1 = 32'd20
; 
32'd8013: dataIn1 = 32'd23
; 
32'd8014: dataIn1 = 32'd24
; 
32'd8015: dataIn1 = 32'd25
; 
32'd8016: dataIn1 = 32'd27
; 
32'd8017: dataIn1 = 32'd29
; 
32'd8018: dataIn1 = 32'd31
; 
32'd8019: dataIn1 = 32'd1
; 
32'd8020: dataIn1 = 32'd2
; 
32'd8021: dataIn1 = 32'd3
; 
32'd8022: dataIn1 = 32'd4
; 
32'd8023: dataIn1 = 32'd5
; 
32'd8024: dataIn1 = 32'd6
; 
32'd8025: dataIn1 = 32'd8
; 
32'd8026: dataIn1 = 32'd11
; 
32'd8027: dataIn1 = 32'd12
; 
32'd8028: dataIn1 = 32'd13
; 
32'd8029: dataIn1 = 32'd18
; 
32'd8030: dataIn1 = 32'd19
; 
32'd8031: dataIn1 = 32'd20
; 
32'd8032: dataIn1 = 32'd21
; 
32'd8033: dataIn1 = 32'd23
; 
32'd8034: dataIn1 = 32'd24
; 
32'd8035: dataIn1 = 32'd25
; 
32'd8036: dataIn1 = 32'd26
; 
32'd8037: dataIn1 = 32'd30
; 
32'd8038: dataIn1 = 32'd31
; 
32'd8039: dataIn1 = 32'd0
; 
32'd8040: dataIn1 = 32'd1
; 
32'd8041: dataIn1 = 32'd3
; 
32'd8042: dataIn1 = 32'd6
; 
32'd8043: dataIn1 = 32'd7
; 
32'd8044: dataIn1 = 32'd9
; 
32'd8045: dataIn1 = 32'd11
; 
32'd8046: dataIn1 = 32'd12
; 
32'd8047: dataIn1 = 32'd13
; 
32'd8048: dataIn1 = 32'd14
; 
32'd8049: dataIn1 = 32'd15
; 
32'd8050: dataIn1 = 32'd17
; 
32'd8051: dataIn1 = 32'd20
; 
32'd8052: dataIn1 = 32'd22
; 
32'd8053: dataIn1 = 32'd23
; 
32'd8054: dataIn1 = 32'd24
; 
32'd8055: dataIn1 = 32'd26
; 
32'd8056: dataIn1 = 32'd27
; 
32'd8057: dataIn1 = 32'd31
; 
32'd8058: dataIn1 = 32'd0
; 
32'd8059: dataIn1 = 32'd1
; 
32'd8060: dataIn1 = 32'd2
; 
32'd8061: dataIn1 = 32'd3
; 
32'd8062: dataIn1 = 32'd4
; 
32'd8063: dataIn1 = 32'd5
; 
32'd8064: dataIn1 = 32'd7
; 
32'd8065: dataIn1 = 32'd11
; 
32'd8066: dataIn1 = 32'd12
; 
32'd8067: dataIn1 = 32'd15
; 
32'd8068: dataIn1 = 32'd18
; 
32'd8069: dataIn1 = 32'd19
; 
32'd8070: dataIn1 = 32'd20
; 
32'd8071: dataIn1 = 32'd21
; 
32'd8072: dataIn1 = 32'd22
; 
32'd8073: dataIn1 = 32'd23
; 
32'd8074: dataIn1 = 32'd24
; 
32'd8075: dataIn1 = 32'd25
; 
32'd8076: dataIn1 = 32'd26
; 
32'd8077: dataIn1 = 32'd28
; 
32'd8078: dataIn1 = 32'd29
; 
32'd8079: dataIn1 = 32'd1
; 
32'd8080: dataIn1 = 32'd2
; 
32'd8081: dataIn1 = 32'd3
; 
32'd8082: dataIn1 = 32'd4
; 
32'd8083: dataIn1 = 32'd5
; 
32'd8084: dataIn1 = 32'd7
; 
32'd8085: dataIn1 = 32'd8
; 
32'd8086: dataIn1 = 32'd10
; 
32'd8087: dataIn1 = 32'd11
; 
32'd8088: dataIn1 = 32'd12
; 
32'd8089: dataIn1 = 32'd13
; 
32'd8090: dataIn1 = 32'd14
; 
32'd8091: dataIn1 = 32'd16
; 
32'd8092: dataIn1 = 32'd17
; 
32'd8093: dataIn1 = 32'd18
; 
32'd8094: dataIn1 = 32'd19
; 
32'd8095: dataIn1 = 32'd21
; 
32'd8096: dataIn1 = 32'd23
; 
32'd8097: dataIn1 = 32'd24
; 
32'd8098: dataIn1 = 32'd25
; 
32'd8099: dataIn1 = 32'd26
; 
32'd8100: dataIn1 = 32'd27
; 
32'd8101: dataIn1 = 32'd28
; 
32'd8102: dataIn1 = 32'd29
; 
32'd8103: dataIn1 = 32'd31
; 
32'd8104: dataIn1 = 32'd1
; 
32'd8105: dataIn1 = 32'd2
; 
32'd8106: dataIn1 = 32'd5
; 
32'd8107: dataIn1 = 32'd6
; 
32'd8108: dataIn1 = 32'd12
; 
32'd8109: dataIn1 = 32'd13
; 
32'd8110: dataIn1 = 32'd15
; 
32'd8111: dataIn1 = 32'd16
; 
32'd8112: dataIn1 = 32'd20
; 
32'd8113: dataIn1 = 32'd21
; 
32'd8114: dataIn1 = 32'd23
; 
32'd8115: dataIn1 = 32'd24
; 
32'd8116: dataIn1 = 32'd26
; 
32'd8117: dataIn1 = 32'd27
; 
32'd8118: dataIn1 = 32'd29
; 
32'd8119: dataIn1 = 32'd30
; 
32'd8120: dataIn1 = 32'd31
; 
32'd8121: dataIn1 = 32'd1
; 
32'd8122: dataIn1 = 32'd3
; 
32'd8123: dataIn1 = 32'd4
; 
32'd8124: dataIn1 = 32'd5
; 
32'd8125: dataIn1 = 32'd7
; 
32'd8126: dataIn1 = 32'd8
; 
32'd8127: dataIn1 = 32'd9
; 
32'd8128: dataIn1 = 32'd10
; 
32'd8129: dataIn1 = 32'd11
; 
32'd8130: dataIn1 = 32'd14
; 
32'd8131: dataIn1 = 32'd16
; 
32'd8132: dataIn1 = 32'd17
; 
32'd8133: dataIn1 = 32'd18
; 
32'd8134: dataIn1 = 32'd19
; 
32'd8135: dataIn1 = 32'd21
; 
32'd8136: dataIn1 = 32'd22
; 
32'd8137: dataIn1 = 32'd25
; 
32'd8138: dataIn1 = 32'd27
; 
32'd8139: dataIn1 = 32'd28
; 
32'd8140: dataIn1 = 32'd29
; 
32'd8141: dataIn1 = 32'd30
; 
32'd8142: dataIn1 = 32'd31
; 
32'd8143: dataIn1 = 32'd0
; 
32'd8144: dataIn1 = 32'd2
; 
32'd8145: dataIn1 = 32'd4
; 
32'd8146: dataIn1 = 32'd6
; 
32'd8147: dataIn1 = 32'd8
; 
32'd8148: dataIn1 = 32'd11
; 
32'd8149: dataIn1 = 32'd12
; 
32'd8150: dataIn1 = 32'd13
; 
32'd8151: dataIn1 = 32'd14
; 
32'd8152: dataIn1 = 32'd15
; 
32'd8153: dataIn1 = 32'd18
; 
32'd8154: dataIn1 = 32'd19
; 
32'd8155: dataIn1 = 32'd21
; 
32'd8156: dataIn1 = 32'd22
; 
32'd8157: dataIn1 = 32'd23
; 
32'd8158: dataIn1 = 32'd25
; 
32'd8159: dataIn1 = 32'd26
; 
32'd8160: dataIn1 = 32'd27
; 
32'd8161: dataIn1 = 32'd28
; 
32'd8162: dataIn1 = 32'd29
; 
32'd8163: dataIn1 = 32'd30
; 
32'd8164: dataIn1 = 32'd1
; 
32'd8165: dataIn1 = 32'd4
; 
32'd8166: dataIn1 = 32'd7
; 
32'd8167: dataIn1 = 32'd8
; 
32'd8168: dataIn1 = 32'd9
; 
32'd8169: dataIn1 = 32'd11
; 
32'd8170: dataIn1 = 32'd12
; 
32'd8171: dataIn1 = 32'd15
; 
32'd8172: dataIn1 = 32'd17
; 
32'd8173: dataIn1 = 32'd19
; 
32'd8174: dataIn1 = 32'd20
; 
32'd8175: dataIn1 = 32'd21
; 
32'd8176: dataIn1 = 32'd23
; 
32'd8177: dataIn1 = 32'd24
; 
32'd8178: dataIn1 = 32'd27
; 
32'd8179: dataIn1 = 32'd29
; 
32'd8180: dataIn1 = 32'd30
; 
32'd8181: dataIn1 = 32'd31
; 
32'd8182: dataIn1 = 32'd2
; 
32'd8183: dataIn1 = 32'd3
; 
32'd8184: dataIn1 = 32'd4
; 
32'd8185: dataIn1 = 32'd5
; 
32'd8186: dataIn1 = 32'd7
; 
32'd8187: dataIn1 = 32'd8
; 
32'd8188: dataIn1 = 32'd9
; 
32'd8189: dataIn1 = 32'd11
; 
32'd8190: dataIn1 = 32'd12
; 
32'd8191: dataIn1 = 32'd13
; 
32'd8192: dataIn1 = 32'd15
; 
32'd8193: dataIn1 = 32'd18
; 
32'd8194: dataIn1 = 32'd19
; 
32'd8195: dataIn1 = 32'd20
; 
32'd8196: dataIn1 = 32'd22
; 
32'd8197: dataIn1 = 32'd24
; 
32'd8198: dataIn1 = 32'd27
; 
32'd8199: dataIn1 = 32'd28
; 
32'd8200: dataIn1 = 32'd29
; 
32'd8201: dataIn1 = 32'd30
; 
32'd8202: dataIn1 = 32'd31
; 
32'd8203: dataIn1 = 32'd0
; 
32'd8204: dataIn1 = 32'd1
; 
32'd8205: dataIn1 = 32'd3
; 
32'd8206: dataIn1 = 32'd4
; 
32'd8207: dataIn1 = 32'd6
; 
32'd8208: dataIn1 = 32'd8
; 
32'd8209: dataIn1 = 32'd9
; 
32'd8210: dataIn1 = 32'd10
; 
32'd8211: dataIn1 = 32'd12
; 
32'd8212: dataIn1 = 32'd13
; 
32'd8213: dataIn1 = 32'd14
; 
32'd8214: dataIn1 = 32'd16
; 
32'd8215: dataIn1 = 32'd17
; 
32'd8216: dataIn1 = 32'd18
; 
32'd8217: dataIn1 = 32'd20
; 
32'd8218: dataIn1 = 32'd21
; 
32'd8219: dataIn1 = 32'd24
; 
32'd8220: dataIn1 = 32'd26
; 
32'd8221: dataIn1 = 32'd27
; 
32'd8222: dataIn1 = 32'd28
; 
32'd8223: dataIn1 = 32'd31
; 
32'd8224: dataIn1 = 32'd1
; 
32'd8225: dataIn1 = 32'd2
; 
32'd8226: dataIn1 = 32'd3
; 
32'd8227: dataIn1 = 32'd4
; 
32'd8228: dataIn1 = 32'd6
; 
32'd8229: dataIn1 = 32'd10
; 
32'd8230: dataIn1 = 32'd12
; 
32'd8231: dataIn1 = 32'd16
; 
32'd8232: dataIn1 = 32'd17
; 
32'd8233: dataIn1 = 32'd21
; 
32'd8234: dataIn1 = 32'd23
; 
32'd8235: dataIn1 = 32'd25
; 
32'd8236: dataIn1 = 32'd30
; 
32'd8237: dataIn1 = 32'd1
; 
32'd8238: dataIn1 = 32'd5
; 
32'd8239: dataIn1 = 32'd6
; 
32'd8240: dataIn1 = 32'd7
; 
32'd8241: dataIn1 = 32'd8
; 
32'd8242: dataIn1 = 32'd9
; 
32'd8243: dataIn1 = 32'd10
; 
32'd8244: dataIn1 = 32'd11
; 
32'd8245: dataIn1 = 32'd14
; 
32'd8246: dataIn1 = 32'd19
; 
32'd8247: dataIn1 = 32'd21
; 
32'd8248: dataIn1 = 32'd22
; 
32'd8249: dataIn1 = 32'd23
; 
32'd8250: dataIn1 = 32'd26
; 
32'd8251: dataIn1 = 32'd27
; 
32'd8252: dataIn1 = 32'd29
; 
32'd8253: dataIn1 = 32'd30
; 
32'd8254: dataIn1 = 32'd0
; 
32'd8255: dataIn1 = 32'd3
; 
32'd8256: dataIn1 = 32'd4
; 
32'd8257: dataIn1 = 32'd5
; 
32'd8258: dataIn1 = 32'd6
; 
32'd8259: dataIn1 = 32'd7
; 
32'd8260: dataIn1 = 32'd8
; 
32'd8261: dataIn1 = 32'd9
; 
32'd8262: dataIn1 = 32'd13
; 
32'd8263: dataIn1 = 32'd15
; 
32'd8264: dataIn1 = 32'd18
; 
32'd8265: dataIn1 = 32'd19
; 
32'd8266: dataIn1 = 32'd20
; 
32'd8267: dataIn1 = 32'd21
; 
32'd8268: dataIn1 = 32'd23
; 
32'd8269: dataIn1 = 32'd25
; 
32'd8270: dataIn1 = 32'd28
; 
32'd8271: dataIn1 = 32'd30
; 
32'd8272: dataIn1 = 32'd0
; 
32'd8273: dataIn1 = 32'd2
; 
32'd8274: dataIn1 = 32'd3
; 
32'd8275: dataIn1 = 32'd5
; 
32'd8276: dataIn1 = 32'd8
; 
32'd8277: dataIn1 = 32'd10
; 
32'd8278: dataIn1 = 32'd15
; 
32'd8279: dataIn1 = 32'd16
; 
32'd8280: dataIn1 = 32'd17
; 
32'd8281: dataIn1 = 32'd18
; 
32'd8282: dataIn1 = 32'd19
; 
32'd8283: dataIn1 = 32'd20
; 
32'd8284: dataIn1 = 32'd21
; 
32'd8285: dataIn1 = 32'd22
; 
32'd8286: dataIn1 = 32'd26
; 
32'd8287: dataIn1 = 32'd27
; 
32'd8288: dataIn1 = 32'd28
; 
32'd8289: dataIn1 = 32'd31
; 
32'd8290: dataIn1 = 32'd0
; 
32'd8291: dataIn1 = 32'd1
; 
32'd8292: dataIn1 = 32'd3
; 
32'd8293: dataIn1 = 32'd8
; 
32'd8294: dataIn1 = 32'd9
; 
32'd8295: dataIn1 = 32'd10
; 
32'd8296: dataIn1 = 32'd11
; 
32'd8297: dataIn1 = 32'd12
; 
32'd8298: dataIn1 = 32'd13
; 
32'd8299: dataIn1 = 32'd14
; 
32'd8300: dataIn1 = 32'd22
; 
32'd8301: dataIn1 = 32'd24
; 
32'd8302: dataIn1 = 32'd25
; 
32'd8303: dataIn1 = 32'd28
; 
32'd8304: dataIn1 = 32'd29
; 
32'd8305: dataIn1 = 32'd30
; 
32'd8306: dataIn1 = 32'd31
; 
32'd8307: dataIn1 = 32'd1
; 
32'd8308: dataIn1 = 32'd2
; 
32'd8309: dataIn1 = 32'd4
; 
32'd8310: dataIn1 = 32'd5
; 
32'd8311: dataIn1 = 32'd7
; 
32'd8312: dataIn1 = 32'd9
; 
32'd8313: dataIn1 = 32'd10
; 
32'd8314: dataIn1 = 32'd12
; 
32'd8315: dataIn1 = 32'd13
; 
32'd8316: dataIn1 = 32'd14
; 
32'd8317: dataIn1 = 32'd19
; 
32'd8318: dataIn1 = 32'd20
; 
32'd8319: dataIn1 = 32'd21
; 
32'd8320: dataIn1 = 32'd22
; 
32'd8321: dataIn1 = 32'd23
; 
32'd8322: dataIn1 = 32'd25
; 
32'd8323: dataIn1 = 32'd26
; 
32'd8324: dataIn1 = 32'd29
; 
32'd8325: dataIn1 = 32'd30
; 
32'd8326: dataIn1 = 32'd31
; 
32'd8327: dataIn1 = 32'd0
; 
32'd8328: dataIn1 = 32'd1
; 
32'd8329: dataIn1 = 32'd4
; 
32'd8330: dataIn1 = 32'd5
; 
32'd8331: dataIn1 = 32'd7
; 
32'd8332: dataIn1 = 32'd8
; 
32'd8333: dataIn1 = 32'd12
; 
32'd8334: dataIn1 = 32'd14
; 
32'd8335: dataIn1 = 32'd16
; 
32'd8336: dataIn1 = 32'd17
; 
32'd8337: dataIn1 = 32'd18
; 
32'd8338: dataIn1 = 32'd19
; 
32'd8339: dataIn1 = 32'd23
; 
32'd8340: dataIn1 = 32'd24
; 
32'd8341: dataIn1 = 32'd25
; 
32'd8342: dataIn1 = 32'd26
; 
32'd8343: dataIn1 = 32'd27
; 
32'd8344: dataIn1 = 32'd28
; 
32'd8345: dataIn1 = 32'd29
; 
32'd8346: dataIn1 = 32'd30
; 
32'd8347: dataIn1 = 32'd31
; 
32'd8348: dataIn1 = 32'd0
; 
32'd8349: dataIn1 = 32'd2
; 
32'd8350: dataIn1 = 32'd3
; 
32'd8351: dataIn1 = 32'd6
; 
32'd8352: dataIn1 = 32'd9
; 
32'd8353: dataIn1 = 32'd10
; 
32'd8354: dataIn1 = 32'd11
; 
32'd8355: dataIn1 = 32'd12
; 
32'd8356: dataIn1 = 32'd15
; 
32'd8357: dataIn1 = 32'd17
; 
32'd8358: dataIn1 = 32'd20
; 
32'd8359: dataIn1 = 32'd22
; 
32'd8360: dataIn1 = 32'd23
; 
32'd8361: dataIn1 = 32'd24
; 
32'd8362: dataIn1 = 32'd26
; 
32'd8363: dataIn1 = 32'd27
; 
32'd8364: dataIn1 = 32'd29
; 
32'd8365: dataIn1 = 32'd30
; 
32'd8366: dataIn1 = 32'd31
; 
32'd8367: dataIn1 = 32'd1
; 
32'd8368: dataIn1 = 32'd3
; 
32'd8369: dataIn1 = 32'd4
; 
32'd8370: dataIn1 = 32'd5
; 
32'd8371: dataIn1 = 32'd8
; 
32'd8372: dataIn1 = 32'd12
; 
32'd8373: dataIn1 = 32'd14
; 
32'd8374: dataIn1 = 32'd17
; 
32'd8375: dataIn1 = 32'd18
; 
32'd8376: dataIn1 = 32'd19
; 
32'd8377: dataIn1 = 32'd23
; 
32'd8378: dataIn1 = 32'd27
; 
32'd8379: dataIn1 = 32'd28
; 
32'd8380: dataIn1 = 32'd30
; 
32'd8381: dataIn1 = 32'd31
; 
32'd8382: dataIn1 = 32'd0
; 
32'd8383: dataIn1 = 32'd1
; 
32'd8384: dataIn1 = 32'd3
; 
32'd8385: dataIn1 = 32'd5
; 
32'd8386: dataIn1 = 32'd6
; 
32'd8387: dataIn1 = 32'd7
; 
32'd8388: dataIn1 = 32'd8
; 
32'd8389: dataIn1 = 32'd9
; 
32'd8390: dataIn1 = 32'd10
; 
32'd8391: dataIn1 = 32'd11
; 
32'd8392: dataIn1 = 32'd13
; 
32'd8393: dataIn1 = 32'd14
; 
32'd8394: dataIn1 = 32'd15
; 
32'd8395: dataIn1 = 32'd16
; 
32'd8396: dataIn1 = 32'd17
; 
32'd8397: dataIn1 = 32'd18
; 
32'd8398: dataIn1 = 32'd19
; 
32'd8399: dataIn1 = 32'd20
; 
32'd8400: dataIn1 = 32'd21
; 
32'd8401: dataIn1 = 32'd23
; 
32'd8402: dataIn1 = 32'd25
; 
32'd8403: dataIn1 = 32'd26
; 
32'd8404: dataIn1 = 32'd27
; 
32'd8405: dataIn1 = 32'd31
; 
32'd8406: dataIn1 = 32'd0
; 
32'd8407: dataIn1 = 32'd3
; 
32'd8408: dataIn1 = 32'd4
; 
32'd8409: dataIn1 = 32'd5
; 
32'd8410: dataIn1 = 32'd6
; 
32'd8411: dataIn1 = 32'd7
; 
32'd8412: dataIn1 = 32'd8
; 
32'd8413: dataIn1 = 32'd9
; 
32'd8414: dataIn1 = 32'd12
; 
32'd8415: dataIn1 = 32'd15
; 
32'd8416: dataIn1 = 32'd16
; 
32'd8417: dataIn1 = 32'd17
; 
32'd8418: dataIn1 = 32'd18
; 
32'd8419: dataIn1 = 32'd22
; 
32'd8420: dataIn1 = 32'd25
; 
32'd8421: dataIn1 = 32'd26
; 
32'd8422: dataIn1 = 32'd27
; 
32'd8423: dataIn1 = 32'd28
; 
32'd8424: dataIn1 = 32'd29
; 
32'd8425: dataIn1 = 32'd31
; 
32'd8426: dataIn1 = 32'd1
; 
32'd8427: dataIn1 = 32'd2
; 
32'd8428: dataIn1 = 32'd3
; 
32'd8429: dataIn1 = 32'd4
; 
32'd8430: dataIn1 = 32'd5
; 
32'd8431: dataIn1 = 32'd6
; 
32'd8432: dataIn1 = 32'd10
; 
32'd8433: dataIn1 = 32'd14
; 
32'd8434: dataIn1 = 32'd16
; 
32'd8435: dataIn1 = 32'd17
; 
32'd8436: dataIn1 = 32'd18
; 
32'd8437: dataIn1 = 32'd19
; 
32'd8438: dataIn1 = 32'd20
; 
32'd8439: dataIn1 = 32'd21
; 
32'd8440: dataIn1 = 32'd22
; 
32'd8441: dataIn1 = 32'd24
; 
32'd8442: dataIn1 = 32'd27
; 
32'd8443: dataIn1 = 32'd29
; 
32'd8444: dataIn1 = 32'd30
; 
32'd8445: dataIn1 = 32'd1
; 
32'd8446: dataIn1 = 32'd3
; 
32'd8447: dataIn1 = 32'd4
; 
32'd8448: dataIn1 = 32'd5
; 
32'd8449: dataIn1 = 32'd6
; 
32'd8450: dataIn1 = 32'd9
; 
32'd8451: dataIn1 = 32'd10
; 
32'd8452: dataIn1 = 32'd11
; 
32'd8453: dataIn1 = 32'd16
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd60; 
32'd3: dataIn2 = 32'd85; 
32'd4: dataIn2 = 32'd20; 
32'd5: dataIn2 = 32'd61; 
32'd6: dataIn2 = 32'd47; 
32'd7: dataIn2 = 32'd41; 
32'd8: dataIn2 = 32'd98; 
32'd9: dataIn2 = 32'd85; 
32'd10: dataIn2 = 32'd20; 
32'd11: dataIn2 = 32'd1; 
32'd12: dataIn2 = 32'd59; 
32'd13: dataIn2 = 32'd58; 
32'd14: dataIn2 = 32'd71; 
32'd15: dataIn2 = 32'd63; 
32'd16: dataIn2 = 32'd96; 
32'd17: dataIn2 = 32'd81; 
32'd18: dataIn2 = 32'd85; 
32'd19: dataIn2 = 32'd50; 
32'd20: dataIn2 = 32'd35; 
32'd21: dataIn2 = 32'd60; 
32'd22: dataIn2 = 32'd14; 
32'd23: dataIn2 = 32'd62; 
32'd24: dataIn2 = 32'd62; 
32'd25: dataIn2 = 32'd36; 
32'd26: dataIn2 = 32'd49; 
32'd27: dataIn2 = 32'd51; 
32'd28: dataIn2 = 32'd68; 
32'd29: dataIn2 = 32'd73; 
32'd30: dataIn2 = 32'd52; 
32'd31: dataIn2 = 32'd84; 
32'd32: dataIn2 = 32'd88; 
32'd33: dataIn2 = 32'd20; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd170: dataIn2 = 32'd98; 
32'd171: dataIn2 = 32'd2; 
32'd172: dataIn2 = 32'd19; 
32'd173: dataIn2 = 32'd17; 
32'd174: dataIn2 = 32'd91; 
32'd175: dataIn2 = 32'd53; 
32'd176: dataIn2 = 32'd29; 
32'd177: dataIn2 = 32'd66; 
32'd178: dataIn2 = 32'd85; 
32'd179: dataIn2 = 32'd77; 
32'd180: dataIn2 = 32'd34; 
32'd181: dataIn2 = 32'd42; 
32'd182: dataIn2 = 32'd98; 
32'd183: dataIn2 = 32'd22; 
32'd184: dataIn2 = 32'd37; 
32'd185: dataIn2 = 32'd49; 
32'd186: dataIn2 = 32'd15; 
32'd187: dataIn2 = 32'd20; 
32'd188: dataIn2 = 32'd34; 
32'd189: dataIn2 = 32'd81; 
32'd190: dataIn2 = 32'd96; 
32'd191: dataIn2 = 32'd79; 
32'd192: dataIn2 = 32'd26; 
32'd193: dataIn2 = 32'd90; 
32'd194: dataIn2 = 32'd83; 
32'd195: dataIn2 = 32'd62; 
32'd196: dataIn2 = 32'd59; 
32'd197: dataIn2 = 32'd65; 
32'd198: dataIn2 = 32'd20; 
32'd199: dataIn2 = 32'd7; 
32'd200: dataIn2 = 32'd98; 
32'd201: dataIn2 = 32'd58; 
32'd202: dataIn2 = 32'd11; 
32'd203: dataIn2 = 32'd26; 
32'd204: dataIn2 = 32'd29; 
32'd205: dataIn2 = 32'd86; 
32'd206: dataIn2 = 32'd59; 
32'd207: dataIn2 = 32'd77; 
32'd208: dataIn2 = 32'd21; 
32'd209: dataIn2 = 32'd0; 
32'd210: dataIn2 = 32'd67; 
32'd211: dataIn2 = 32'd92; 
32'd212: dataIn2 = 32'd2; 
32'd213: dataIn2 = 32'd57; 
32'd214: dataIn2 = 32'd43; 
32'd215: dataIn2 = 32'd26; 
32'd216: dataIn2 = 32'd26; 
32'd217: dataIn2 = 32'd50; 
32'd218: dataIn2 = 32'd49; 
32'd219: dataIn2 = 32'd47; 
32'd220: dataIn2 = 32'd41; 
32'd221: dataIn2 = 32'd74; 
32'd222: dataIn2 = 32'd88; 
32'd223: dataIn2 = 32'd17; 
32'd224: dataIn2 = 32'd18; 
32'd225: dataIn2 = 32'd61; 
32'd226: dataIn2 = 32'd65; 
32'd227: dataIn2 = 32'd75; 
32'd228: dataIn2 = 32'd99; 
32'd229: dataIn2 = 32'd18; 
32'd230: dataIn2 = 32'd83; 
32'd231: dataIn2 = 32'd95; 
32'd232: dataIn2 = 32'd16; 
32'd233: dataIn2 = 32'd9; 
32'd234: dataIn2 = 32'd60; 
32'd235: dataIn2 = 32'd62; 
32'd236: dataIn2 = 32'd63; 
32'd237: dataIn2 = 32'd76; 
32'd238: dataIn2 = 32'd63; 
32'd239: dataIn2 = 32'd49; 
32'd240: dataIn2 = 32'd0; 
32'd241: dataIn2 = 32'd76; 
32'd242: dataIn2 = 32'd26; 
32'd243: dataIn2 = 32'd8; 
32'd244: dataIn2 = 32'd4; 
32'd245: dataIn2 = 32'd100; 
32'd246: dataIn2 = 32'd95; 
32'd247: dataIn2 = 32'd56; 
32'd248: dataIn2 = 32'd36; 
32'd249: dataIn2 = 32'd97; 
32'd250: dataIn2 = 32'd70; 
32'd251: dataIn2 = 32'd48; 
32'd252: dataIn2 = 32'd7; 
32'd253: dataIn2 = 32'd2; 
32'd254: dataIn2 = 32'd36; 
32'd255: dataIn2 = 32'd10; 
32'd256: dataIn2 = 32'd68; 
32'd257: dataIn2 = 32'd49; 
32'd258: dataIn2 = 32'd47; 
32'd259: dataIn2 = 32'd54; 
32'd260: dataIn2 = 32'd33; 
32'd261: dataIn2 = 32'd76; 
32'd262: dataIn2 = 32'd10; 
32'd263: dataIn2 = 32'd41; 
32'd264: dataIn2 = 32'd76; 
32'd265: dataIn2 = 32'd55; 
32'd266: dataIn2 = 32'd98; 
32'd267: dataIn2 = 32'd18; 
32'd268: dataIn2 = 32'd96; 
32'd269: dataIn2 = 32'd27; 
32'd270: dataIn2 = 32'd42; 
32'd271: dataIn2 = 32'd75; 
32'd272: dataIn2 = 32'd5; 
32'd273: dataIn2 = 32'd0; 
32'd274: dataIn2 = 32'd48; 
32'd275: dataIn2 = 32'd65; 
32'd276: dataIn2 = 32'd95; 
32'd277: dataIn2 = 32'd84; 
32'd278: dataIn2 = 32'd66; 
32'd279: dataIn2 = 32'd16; 
32'd280: dataIn2 = 32'd28; 
32'd281: dataIn2 = 32'd79; 
32'd282: dataIn2 = 32'd41; 
32'd283: dataIn2 = 32'd94; 
32'd284: dataIn2 = 32'd23; 
32'd285: dataIn2 = 32'd47; 
32'd286: dataIn2 = 32'd73; 
32'd287: dataIn2 = 32'd45; 
32'd288: dataIn2 = 32'd84; 
32'd289: dataIn2 = 32'd16; 
32'd290: dataIn2 = 32'd78; 
32'd291: dataIn2 = 32'd99; 
32'd292: dataIn2 = 32'd75; 
32'd293: dataIn2 = 32'd97; 
32'd294: dataIn2 = 32'd43; 
32'd295: dataIn2 = 32'd65; 
32'd296: dataIn2 = 32'd6; 
32'd297: dataIn2 = 32'd37; 
32'd298: dataIn2 = 32'd31; 
32'd299: dataIn2 = 32'd90; 
32'd300: dataIn2 = 32'd27; 
32'd301: dataIn2 = 32'd62; 
32'd302: dataIn2 = 32'd5; 
32'd303: dataIn2 = 32'd46; 
32'd304: dataIn2 = 32'd37; 
32'd305: dataIn2 = 32'd17; 
32'd306: dataIn2 = 32'd86; 
32'd307: dataIn2 = 32'd58; 
32'd308: dataIn2 = 32'd53; 
32'd309: dataIn2 = 32'd0; 
32'd310: dataIn2 = 32'd50; 
32'd311: dataIn2 = 32'd28; 
32'd312: dataIn2 = 32'd99; 
32'd313: dataIn2 = 32'd29; 
32'd314: dataIn2 = 32'd79; 
32'd315: dataIn2 = 32'd30; 
32'd316: dataIn2 = 32'd72; 
32'd317: dataIn2 = 32'd4; 
32'd318: dataIn2 = 32'd12; 
32'd319: dataIn2 = 32'd73; 
32'd320: dataIn2 = 32'd35; 
32'd321: dataIn2 = 32'd70; 
32'd322: dataIn2 = 32'd92; 
32'd323: dataIn2 = 32'd97; 
32'd324: dataIn2 = 32'd80; 
32'd325: dataIn2 = 32'd50; 
32'd326: dataIn2 = 32'd23; 
32'd327: dataIn2 = 32'd31; 
32'd328: dataIn2 = 32'd48; 
32'd329: dataIn2 = 32'd86; 
32'd330: dataIn2 = 32'd2; 
32'd331: dataIn2 = 32'd84; 
32'd332: dataIn2 = 32'd23; 
32'd333: dataIn2 = 32'd87; 
32'd334: dataIn2 = 32'd7; 
32'd335: dataIn2 = 32'd97; 
32'd336: dataIn2 = 32'd5; 
32'd337: dataIn2 = 32'd22; 
32'd338: dataIn2 = 32'd72; 
32'd339: dataIn2 = 32'd79; 
32'd340: dataIn2 = 32'd46; 
32'd341: dataIn2 = 32'd85; 
32'd342: dataIn2 = 32'd5; 
32'd343: dataIn2 = 32'd22; 
32'd344: dataIn2 = 32'd99; 
32'd345: dataIn2 = 32'd90; 
32'd346: dataIn2 = 32'd26; 
32'd347: dataIn2 = 32'd63; 
32'd348: dataIn2 = 32'd58; 
32'd349: dataIn2 = 32'd95; 
32'd350: dataIn2 = 32'd100; 
32'd351: dataIn2 = 32'd60; 
32'd352: dataIn2 = 32'd99; 
32'd353: dataIn2 = 32'd13; 
32'd354: dataIn2 = 32'd6; 
32'd355: dataIn2 = 32'd79; 
32'd356: dataIn2 = 32'd49; 
32'd357: dataIn2 = 32'd20; 
32'd358: dataIn2 = 32'd29; 
32'd359: dataIn2 = 32'd52; 
32'd360: dataIn2 = 32'd86; 
32'd361: dataIn2 = 32'd48; 
32'd362: dataIn2 = 32'd36; 
32'd363: dataIn2 = 32'd2; 
32'd364: dataIn2 = 32'd28; 
32'd365: dataIn2 = 32'd64; 
32'd366: dataIn2 = 32'd20; 
32'd367: dataIn2 = 32'd31; 
32'd368: dataIn2 = 32'd74; 
32'd369: dataIn2 = 32'd80; 
32'd370: dataIn2 = 32'd65; 
32'd371: dataIn2 = 32'd78; 
32'd372: dataIn2 = 32'd97; 
32'd373: dataIn2 = 32'd95; 
32'd374: dataIn2 = 32'd100; 
32'd375: dataIn2 = 32'd78; 
32'd376: dataIn2 = 32'd73; 
32'd377: dataIn2 = 32'd86; 
32'd378: dataIn2 = 32'd18; 
32'd379: dataIn2 = 32'd1; 
32'd380: dataIn2 = 32'd25; 
32'd381: dataIn2 = 32'd53; 
32'd382: dataIn2 = 32'd50; 
32'd383: dataIn2 = 32'd14; 
32'd384: dataIn2 = 32'd3; 
32'd385: dataIn2 = 32'd99; 
32'd386: dataIn2 = 32'd76; 
32'd387: dataIn2 = 32'd40; 
32'd388: dataIn2 = 32'd18; 
32'd389: dataIn2 = 32'd19; 
32'd390: dataIn2 = 32'd49; 
32'd391: dataIn2 = 32'd10; 
32'd392: dataIn2 = 32'd45; 
32'd393: dataIn2 = 32'd97; 
32'd394: dataIn2 = 32'd32; 
32'd395: dataIn2 = 32'd56; 
32'd396: dataIn2 = 32'd64; 
32'd397: dataIn2 = 32'd76; 
32'd398: dataIn2 = 32'd98; 
32'd399: dataIn2 = 32'd15; 
32'd400: dataIn2 = 32'd77; 
32'd401: dataIn2 = 32'd100; 
32'd402: dataIn2 = 32'd87; 
32'd403: dataIn2 = 32'd74; 
32'd404: dataIn2 = 32'd36; 
32'd405: dataIn2 = 32'd43; 
32'd406: dataIn2 = 32'd85; 
32'd407: dataIn2 = 32'd35; 
32'd408: dataIn2 = 32'd55; 
32'd409: dataIn2 = 32'd71; 
32'd410: dataIn2 = 32'd3; 
32'd411: dataIn2 = 32'd57; 
32'd412: dataIn2 = 32'd93; 
32'd413: dataIn2 = 32'd37; 
32'd414: dataIn2 = 32'd98; 
32'd415: dataIn2 = 32'd28; 
32'd416: dataIn2 = 32'd57; 
32'd417: dataIn2 = 32'd60; 
32'd418: dataIn2 = 32'd0; 
32'd419: dataIn2 = 32'd58; 
32'd420: dataIn2 = 32'd33; 
32'd421: dataIn2 = 32'd35; 
32'd422: dataIn2 = 32'd42; 
32'd423: dataIn2 = 32'd18; 
32'd424: dataIn2 = 32'd32; 
32'd425: dataIn2 = 32'd23; 
32'd426: dataIn2 = 32'd62; 
32'd427: dataIn2 = 32'd0; 
32'd428: dataIn2 = 32'd4; 
32'd429: dataIn2 = 32'd21; 
32'd430: dataIn2 = 32'd1; 
32'd431: dataIn2 = 32'd83; 
32'd432: dataIn2 = 32'd96; 
32'd433: dataIn2 = 32'd20; 
32'd434: dataIn2 = 32'd14; 
32'd435: dataIn2 = 32'd36; 
32'd436: dataIn2 = 32'd51; 
32'd437: dataIn2 = 32'd27; 
32'd438: dataIn2 = 32'd29; 
32'd439: dataIn2 = 32'd22; 
32'd440: dataIn2 = 32'd57; 
32'd441: dataIn2 = 32'd30; 
32'd442: dataIn2 = 32'd77; 
32'd443: dataIn2 = 32'd78; 
32'd444: dataIn2 = 32'd82; 
32'd445: dataIn2 = 32'd84; 
32'd446: dataIn2 = 32'd95; 
32'd447: dataIn2 = 32'd27; 
32'd448: dataIn2 = 32'd78; 
32'd449: dataIn2 = 32'd72; 
32'd450: dataIn2 = 32'd96; 
32'd451: dataIn2 = 32'd50; 
32'd452: dataIn2 = 32'd78; 
32'd453: dataIn2 = 32'd88; 
32'd454: dataIn2 = 32'd7; 
32'd455: dataIn2 = 32'd71; 
32'd456: dataIn2 = 32'd38; 
32'd457: dataIn2 = 32'd65; 
32'd458: dataIn2 = 32'd49; 
32'd459: dataIn2 = 32'd21; 
32'd460: dataIn2 = 32'd18; 
32'd461: dataIn2 = 32'd51; 
32'd462: dataIn2 = 32'd52; 
32'd463: dataIn2 = 32'd25; 
32'd464: dataIn2 = 32'd60; 
32'd465: dataIn2 = 32'd69; 
32'd466: dataIn2 = 32'd1; 
32'd467: dataIn2 = 32'd26; 
32'd468: dataIn2 = 32'd12; 
32'd469: dataIn2 = 32'd25; 
32'd470: dataIn2 = 32'd99; 
32'd471: dataIn2 = 32'd37; 
32'd472: dataIn2 = 32'd15; 
32'd473: dataIn2 = 32'd11; 
32'd474: dataIn2 = 32'd24; 
32'd475: dataIn2 = 32'd70; 
32'd476: dataIn2 = 32'd7; 
32'd477: dataIn2 = 32'd7; 
32'd478: dataIn2 = 32'd73; 
32'd479: dataIn2 = 32'd61; 
32'd480: dataIn2 = 32'd58; 
32'd481: dataIn2 = 32'd78; 
32'd482: dataIn2 = 32'd72; 
32'd483: dataIn2 = 32'd51; 
32'd484: dataIn2 = 32'd27; 
32'd485: dataIn2 = 32'd47; 
32'd486: dataIn2 = 32'd50; 
32'd487: dataIn2 = 32'd17; 
32'd488: dataIn2 = 32'd61; 
32'd489: dataIn2 = 32'd68; 
32'd490: dataIn2 = 32'd93; 
32'd491: dataIn2 = 32'd41; 
32'd492: dataIn2 = 32'd18; 
32'd493: dataIn2 = 32'd60; 
32'd494: dataIn2 = 32'd42; 
32'd495: dataIn2 = 32'd81; 
32'd496: dataIn2 = 32'd83; 
32'd497: dataIn2 = 32'd22; 
32'd498: dataIn2 = 32'd35; 
32'd499: dataIn2 = 32'd77; 
32'd500: dataIn2 = 32'd56; 
32'd501: dataIn2 = 32'd67; 
32'd502: dataIn2 = 32'd48; 
32'd503: dataIn2 = 32'd51; 
32'd504: dataIn2 = 32'd42; 
32'd505: dataIn2 = 32'd15; 
32'd506: dataIn2 = 32'd24; 
32'd507: dataIn2 = 32'd100; 
32'd508: dataIn2 = 32'd100; 
32'd509: dataIn2 = 32'd45; 
32'd510: dataIn2 = 32'd79; 
32'd511: dataIn2 = 32'd7; 
32'd512: dataIn2 = 32'd93; 
32'd513: dataIn2 = 32'd93; 
32'd514: dataIn2 = 32'd91; 
32'd515: dataIn2 = 32'd79; 
32'd516: dataIn2 = 32'd75; 
32'd517: dataIn2 = 32'd24; 
32'd518: dataIn2 = 32'd31; 
32'd519: dataIn2 = 32'd38; 
32'd520: dataIn2 = 32'd47; 
32'd521: dataIn2 = 32'd41; 
32'd522: dataIn2 = 32'd96; 
32'd523: dataIn2 = 32'd10; 
32'd524: dataIn2 = 32'd49; 
32'd525: dataIn2 = 32'd99; 
32'd526: dataIn2 = 32'd11; 
32'd527: dataIn2 = 32'd23; 
32'd528: dataIn2 = 32'd7; 
32'd529: dataIn2 = 32'd28; 
32'd530: dataIn2 = 32'd73; 
32'd531: dataIn2 = 32'd48; 
32'd532: dataIn2 = 32'd71; 
32'd533: dataIn2 = 32'd93; 
32'd534: dataIn2 = 32'd54; 
32'd535: dataIn2 = 32'd20; 
32'd536: dataIn2 = 32'd38; 
32'd537: dataIn2 = 32'd8; 
32'd538: dataIn2 = 32'd1; 
32'd539: dataIn2 = 32'd76; 
32'd540: dataIn2 = 32'd53; 
32'd541: dataIn2 = 32'd88; 
32'd542: dataIn2 = 32'd53; 
32'd543: dataIn2 = 32'd58; 
32'd544: dataIn2 = 32'd15; 
32'd545: dataIn2 = 32'd46; 
32'd546: dataIn2 = 32'd38; 
32'd547: dataIn2 = 32'd11; 
32'd548: dataIn2 = 32'd70; 
32'd549: dataIn2 = 32'd88; 
32'd550: dataIn2 = 32'd80; 
32'd551: dataIn2 = 32'd14; 
32'd552: dataIn2 = 32'd44; 
32'd553: dataIn2 = 32'd14; 
32'd554: dataIn2 = 32'd44; 
32'd555: dataIn2 = 32'd7; 
32'd556: dataIn2 = 32'd19; 
32'd557: dataIn2 = 32'd61; 
32'd558: dataIn2 = 32'd94; 
32'd559: dataIn2 = 32'd34; 
32'd560: dataIn2 = 32'd33; 
32'd561: dataIn2 = 32'd42; 
32'd562: dataIn2 = 32'd11; 
32'd563: dataIn2 = 32'd5; 
32'd564: dataIn2 = 32'd98; 
32'd565: dataIn2 = 32'd68; 
32'd566: dataIn2 = 32'd54; 
32'd567: dataIn2 = 32'd36; 
32'd568: dataIn2 = 32'd67; 
32'd569: dataIn2 = 32'd15; 
32'd570: dataIn2 = 32'd2; 
32'd571: dataIn2 = 32'd72; 
32'd572: dataIn2 = 32'd89; 
32'd573: dataIn2 = 32'd51; 
32'd574: dataIn2 = 32'd50; 
32'd575: dataIn2 = 32'd28; 
32'd576: dataIn2 = 32'd76; 
32'd577: dataIn2 = 32'd72; 
32'd578: dataIn2 = 32'd22; 
32'd579: dataIn2 = 32'd40; 
32'd580: dataIn2 = 32'd57; 
32'd581: dataIn2 = 32'd54; 
32'd582: dataIn2 = 32'd2; 
32'd583: dataIn2 = 32'd71; 
32'd584: dataIn2 = 32'd87; 
32'd585: dataIn2 = 32'd28; 
32'd586: dataIn2 = 32'd16; 
32'd587: dataIn2 = 32'd59; 
32'd588: dataIn2 = 32'd73; 
32'd589: dataIn2 = 32'd53; 
32'd590: dataIn2 = 32'd31; 
32'd591: dataIn2 = 32'd87; 
32'd592: dataIn2 = 32'd37; 
32'd593: dataIn2 = 32'd80; 
32'd594: dataIn2 = 32'd42; 
32'd595: dataIn2 = 32'd90; 
32'd596: dataIn2 = 32'd92; 
32'd597: dataIn2 = 32'd81; 
32'd598: dataIn2 = 32'd26; 
32'd599: dataIn2 = 32'd13; 
32'd600: dataIn2 = 32'd88; 
32'd601: dataIn2 = 32'd40; 
32'd602: dataIn2 = 32'd80; 
32'd603: dataIn2 = 32'd21; 
32'd604: dataIn2 = 32'd86; 
32'd605: dataIn2 = 32'd35; 
32'd606: dataIn2 = 32'd38; 
32'd607: dataIn2 = 32'd59; 
32'd608: dataIn2 = 32'd30; 
32'd609: dataIn2 = 32'd45; 
32'd610: dataIn2 = 32'd90; 
32'd611: dataIn2 = 32'd84; 
32'd612: dataIn2 = 32'd35; 
32'd613: dataIn2 = 32'd96; 
32'd614: dataIn2 = 32'd33; 
32'd615: dataIn2 = 32'd72; 
32'd616: dataIn2 = 32'd65; 
32'd617: dataIn2 = 32'd98; 
32'd618: dataIn2 = 32'd64; 
32'd619: dataIn2 = 32'd14; 
32'd620: dataIn2 = 32'd12; 
32'd621: dataIn2 = 32'd73; 
32'd622: dataIn2 = 32'd39; 
32'd623: dataIn2 = 32'd3; 
32'd624: dataIn2 = 32'd57; 
32'd625: dataIn2 = 32'd65; 
32'd626: dataIn2 = 32'd14; 
32'd627: dataIn2 = 32'd43; 
32'd628: dataIn2 = 32'd40; 
32'd629: dataIn2 = 32'd1; 
32'd630: dataIn2 = 32'd22; 
32'd631: dataIn2 = 32'd90; 
32'd632: dataIn2 = 32'd75; 
32'd633: dataIn2 = 32'd54; 
32'd634: dataIn2 = 32'd49; 
32'd635: dataIn2 = 32'd73; 
32'd636: dataIn2 = 32'd47; 
32'd637: dataIn2 = 32'd55; 
32'd638: dataIn2 = 32'd87; 
32'd639: dataIn2 = 32'd13; 
32'd640: dataIn2 = 32'd92; 
32'd641: dataIn2 = 32'd48; 
32'd642: dataIn2 = 32'd1; 
32'd643: dataIn2 = 32'd100; 
32'd644: dataIn2 = 32'd86; 
32'd645: dataIn2 = 32'd2; 
32'd646: dataIn2 = 32'd33; 
32'd647: dataIn2 = 32'd23; 
32'd648: dataIn2 = 32'd6; 
32'd649: dataIn2 = 32'd68; 
32'd650: dataIn2 = 32'd41; 
32'd651: dataIn2 = 32'd35; 
32'd652: dataIn2 = 32'd19; 
32'd653: dataIn2 = 32'd98; 
32'd654: dataIn2 = 32'd77; 
32'd655: dataIn2 = 32'd48; 
32'd656: dataIn2 = 32'd11; 
32'd657: dataIn2 = 32'd88; 
32'd658: dataIn2 = 32'd95; 
32'd659: dataIn2 = 32'd76; 
32'd660: dataIn2 = 32'd24; 
32'd661: dataIn2 = 32'd71; 
32'd662: dataIn2 = 32'd59; 
32'd663: dataIn2 = 32'd22; 
32'd664: dataIn2 = 32'd37; 
32'd665: dataIn2 = 32'd60; 
32'd666: dataIn2 = 32'd36; 
32'd667: dataIn2 = 32'd14; 
32'd668: dataIn2 = 32'd3; 
32'd669: dataIn2 = 32'd23; 
32'd670: dataIn2 = 32'd81; 
32'd671: dataIn2 = 32'd98; 
32'd672: dataIn2 = 32'd0; 
32'd673: dataIn2 = 32'd98; 
32'd674: dataIn2 = 32'd92; 
32'd675: dataIn2 = 32'd55; 
32'd676: dataIn2 = 32'd73; 
32'd677: dataIn2 = 32'd40; 
32'd678: dataIn2 = 32'd23; 
32'd679: dataIn2 = 32'd5; 
32'd680: dataIn2 = 32'd32; 
32'd681: dataIn2 = 32'd40; 
32'd682: dataIn2 = 32'd9; 
32'd683: dataIn2 = 32'd24; 
32'd684: dataIn2 = 32'd62; 
32'd685: dataIn2 = 32'd94; 
32'd686: dataIn2 = 32'd14; 
32'd687: dataIn2 = 32'd3; 
32'd688: dataIn2 = 32'd24; 
32'd689: dataIn2 = 32'd17; 
32'd690: dataIn2 = 32'd70; 
32'd691: dataIn2 = 32'd13; 
32'd692: dataIn2 = 32'd20; 
32'd693: dataIn2 = 32'd13; 
32'd694: dataIn2 = 32'd17; 
32'd695: dataIn2 = 32'd100; 
32'd696: dataIn2 = 32'd51; 
32'd697: dataIn2 = 32'd66; 
32'd698: dataIn2 = 32'd88; 
32'd699: dataIn2 = 32'd94; 
32'd700: dataIn2 = 32'd32; 
32'd701: dataIn2 = 32'd4; 
32'd702: dataIn2 = 32'd55; 
32'd703: dataIn2 = 32'd63; 
32'd704: dataIn2 = 32'd98; 
32'd705: dataIn2 = 32'd11; 
32'd706: dataIn2 = 32'd20; 
32'd707: dataIn2 = 32'd75; 
32'd708: dataIn2 = 32'd19; 
32'd709: dataIn2 = 32'd47; 
32'd710: dataIn2 = 32'd91; 
32'd711: dataIn2 = 32'd14; 
32'd712: dataIn2 = 32'd40; 
32'd713: dataIn2 = 32'd65; 
32'd714: dataIn2 = 32'd87; 
32'd715: dataIn2 = 32'd84; 
32'd716: dataIn2 = 32'd45; 
32'd717: dataIn2 = 32'd70; 
32'd718: dataIn2 = 32'd18; 
32'd719: dataIn2 = 32'd81; 
32'd720: dataIn2 = 32'd87; 
32'd721: dataIn2 = 32'd30; 
32'd722: dataIn2 = 32'd88; 
32'd723: dataIn2 = 32'd26; 
32'd724: dataIn2 = 32'd28; 
32'd725: dataIn2 = 32'd78; 
32'd726: dataIn2 = 32'd15; 
32'd727: dataIn2 = 32'd49; 
32'd728: dataIn2 = 32'd27; 
32'd729: dataIn2 = 32'd94; 
32'd730: dataIn2 = 32'd46; 
32'd731: dataIn2 = 32'd66; 
32'd732: dataIn2 = 32'd75; 
32'd733: dataIn2 = 32'd87; 
32'd734: dataIn2 = 32'd98; 
32'd735: dataIn2 = 32'd82; 
32'd736: dataIn2 = 32'd51; 
32'd737: dataIn2 = 32'd85; 
32'd738: dataIn2 = 32'd56; 
32'd739: dataIn2 = 32'd27; 
32'd740: dataIn2 = 32'd15; 
32'd741: dataIn2 = 32'd32; 
32'd742: dataIn2 = 32'd20; 
32'd743: dataIn2 = 32'd74; 
32'd744: dataIn2 = 32'd89; 
32'd745: dataIn2 = 32'd7; 
32'd746: dataIn2 = 32'd86; 
32'd747: dataIn2 = 32'd82; 
32'd748: dataIn2 = 32'd39; 
32'd749: dataIn2 = 32'd41; 
32'd750: dataIn2 = 32'd51; 
32'd751: dataIn2 = 32'd53; 
32'd752: dataIn2 = 32'd17; 
32'd753: dataIn2 = 32'd62; 
32'd754: dataIn2 = 32'd2; 
32'd755: dataIn2 = 32'd4; 
32'd756: dataIn2 = 32'd87; 
32'd757: dataIn2 = 32'd10; 
32'd758: dataIn2 = 32'd41; 
32'd759: dataIn2 = 32'd29; 
32'd760: dataIn2 = 32'd64; 
32'd761: dataIn2 = 32'd0; 
32'd762: dataIn2 = 32'd48; 
32'd763: dataIn2 = 32'd74; 
32'd764: dataIn2 = 32'd47; 
32'd765: dataIn2 = 32'd55; 
32'd766: dataIn2 = 32'd66; 
32'd767: dataIn2 = 32'd1; 
32'd768: dataIn2 = 32'd82; 
32'd769: dataIn2 = 32'd65; 
32'd770: dataIn2 = 32'd53; 
32'd771: dataIn2 = 32'd2; 
32'd772: dataIn2 = 32'd10; 
32'd773: dataIn2 = 32'd12; 
32'd774: dataIn2 = 32'd38; 
32'd775: dataIn2 = 32'd21; 
32'd776: dataIn2 = 32'd90; 
32'd777: dataIn2 = 32'd33; 
32'd778: dataIn2 = 32'd53; 
32'd779: dataIn2 = 32'd69; 
32'd780: dataIn2 = 32'd75; 
32'd781: dataIn2 = 32'd13; 
32'd782: dataIn2 = 32'd28; 
32'd783: dataIn2 = 32'd35; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_32_40.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
