//64x64 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 2048 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd330 ; 
  wdata_col_base = 32'd23780 ; 
  row_base = 32'd258280 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #220000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd258280: dataIn1 = 32'd0
; 
32'd258281: dataIn1 = 32'd30
; 
32'd258282: dataIn1 = 32'd56
; 
32'd258283: dataIn1 = 32'd90
; 
32'd258284: dataIn1 = 32'd119
; 
32'd258285: dataIn1 = 32'd152
; 
32'd258286: dataIn1 = 32'd178
; 
32'd258287: dataIn1 = 32'd204
; 
32'd258288: dataIn1 = 32'd241
; 
32'd258289: dataIn1 = 32'd278
; 
32'd258290: dataIn1 = 32'd306
; 
32'd258291: dataIn1 = 32'd331
; 
32'd258292: dataIn1 = 32'd360
; 
32'd258293: dataIn1 = 32'd390
; 
32'd258294: dataIn1 = 32'd420
; 
32'd258295: dataIn1 = 32'd451
; 
32'd258296: dataIn1 = 32'd479
; 
32'd258297: dataIn1 = 32'd509
; 
32'd258298: dataIn1 = 32'd535
; 
32'd258299: dataIn1 = 32'd561
; 
32'd258300: dataIn1 = 32'd587
; 
32'd258301: dataIn1 = 32'd620
; 
32'd258302: dataIn1 = 32'd652
; 
32'd258303: dataIn1 = 32'd688
; 
32'd258304: dataIn1 = 32'd714
; 
32'd258305: dataIn1 = 32'd741
; 
32'd258306: dataIn1 = 32'd773
; 
32'd258307: dataIn1 = 32'd804
; 
32'd258308: dataIn1 = 32'd832
; 
32'd258309: dataIn1 = 32'd858
; 
32'd258310: dataIn1 = 32'd890
; 
32'd258311: dataIn1 = 32'd921
; 
32'd258312: dataIn1 = 32'd946
; 
32'd258313: dataIn1 = 32'd977
; 
32'd258314: dataIn1 = 32'd1010
; 
32'd258315: dataIn1 = 32'd1036
; 
32'd258316: dataIn1 = 32'd1063
; 
32'd258317: dataIn1 = 32'd1096
; 
32'd258318: dataIn1 = 32'd1133
; 
32'd258319: dataIn1 = 32'd1167
; 
32'd258320: dataIn1 = 32'd1195
; 
32'd258321: dataIn1 = 32'd1232
; 
32'd258322: dataIn1 = 32'd1264
; 
32'd258323: dataIn1 = 32'd1293
; 
32'd258324: dataIn1 = 32'd1326
; 
32'd258325: dataIn1 = 32'd1356
; 
32'd258326: dataIn1 = 32'd1388
; 
32'd258327: dataIn1 = 32'd1417
; 
32'd258328: dataIn1 = 32'd1445
; 
32'd258329: dataIn1 = 32'd1478
; 
32'd258330: dataIn1 = 32'd1509
; 
32'd258331: dataIn1 = 32'd1544
; 
32'd258332: dataIn1 = 32'd1575
; 
32'd258333: dataIn1 = 32'd1606
; 
32'd258334: dataIn1 = 32'd1639
; 
32'd258335: dataIn1 = 32'd1672
; 
32'd258336: dataIn1 = 32'd1703
; 
32'd258337: dataIn1 = 32'd1735
; 
32'd258338: dataIn1 = 32'd1761
; 
32'd258339: dataIn1 = 32'd1800
; 
32'd258340: dataIn1 = 32'd1835
; 
32'd258341: dataIn1 = 32'd1869
; 
32'd258342: dataIn1 = 32'd1902
; 
32'd258343: dataIn1 = 32'd1934
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd23780: dataIn1 = 32'd0
; 
32'd23781: dataIn1 = 32'd30
; 
32'd23782: dataIn1 = 32'd56
; 
32'd23783: dataIn1 = 32'd90
; 
32'd23784: dataIn1 = 32'd119
; 
32'd23785: dataIn1 = 32'd152
; 
32'd23786: dataIn1 = 32'd178
; 
32'd23787: dataIn1 = 32'd204
; 
32'd23788: dataIn1 = 32'd241
; 
32'd23789: dataIn1 = 32'd278
; 
32'd23790: dataIn1 = 32'd306
; 
32'd23791: dataIn1 = 32'd331
; 
32'd23792: dataIn1 = 32'd360
; 
32'd23793: dataIn1 = 32'd390
; 
32'd23794: dataIn1 = 32'd420
; 
32'd23795: dataIn1 = 32'd451
; 
32'd23796: dataIn1 = 32'd479
; 
32'd23797: dataIn1 = 32'd509
; 
32'd23798: dataIn1 = 32'd535
; 
32'd23799: dataIn1 = 32'd561
; 
32'd23800: dataIn1 = 32'd587
; 
32'd23801: dataIn1 = 32'd620
; 
32'd23802: dataIn1 = 32'd652
; 
32'd23803: dataIn1 = 32'd688
; 
32'd23804: dataIn1 = 32'd714
; 
32'd23805: dataIn1 = 32'd741
; 
32'd23806: dataIn1 = 32'd773
; 
32'd23807: dataIn1 = 32'd804
; 
32'd23808: dataIn1 = 32'd832
; 
32'd23809: dataIn1 = 32'd858
; 
32'd23810: dataIn1 = 32'd890
; 
32'd23811: dataIn1 = 32'd921
; 
32'd23812: dataIn1 = 32'd946
; 
32'd23813: dataIn1 = 32'd977
; 
32'd23814: dataIn1 = 32'd1010
; 
32'd23815: dataIn1 = 32'd1036
; 
32'd23816: dataIn1 = 32'd1063
; 
32'd23817: dataIn1 = 32'd1096
; 
32'd23818: dataIn1 = 32'd1133
; 
32'd23819: dataIn1 = 32'd1167
; 
32'd23820: dataIn1 = 32'd1195
; 
32'd23821: dataIn1 = 32'd1232
; 
32'd23822: dataIn1 = 32'd1264
; 
32'd23823: dataIn1 = 32'd1293
; 
32'd23824: dataIn1 = 32'd1326
; 
32'd23825: dataIn1 = 32'd1356
; 
32'd23826: dataIn1 = 32'd1388
; 
32'd23827: dataIn1 = 32'd1417
; 
32'd23828: dataIn1 = 32'd1445
; 
32'd23829: dataIn1 = 32'd1478
; 
32'd23830: dataIn1 = 32'd1509
; 
32'd23831: dataIn1 = 32'd1544
; 
32'd23832: dataIn1 = 32'd1575
; 
32'd23833: dataIn1 = 32'd1606
; 
32'd23834: dataIn1 = 32'd1639
; 
32'd23835: dataIn1 = 32'd1672
; 
32'd23836: dataIn1 = 32'd1703
; 
32'd23837: dataIn1 = 32'd1735
; 
32'd23838: dataIn1 = 32'd1761
; 
32'd23839: dataIn1 = 32'd1800
; 
32'd23840: dataIn1 = 32'd1835
; 
32'd23841: dataIn1 = 32'd1869
; 
32'd23842: dataIn1 = 32'd1902
; 
32'd23843: dataIn1 = 32'd1934
; 
32'd23844: dataIn1 = 32'd1961
; 
32'd23845: dataIn1 = 32'd1
; 
32'd23846: dataIn1 = 32'd3
; 
32'd23847: dataIn1 = 32'd4
; 
32'd23848: dataIn1 = 32'd7
; 
32'd23849: dataIn1 = 32'd8
; 
32'd23850: dataIn1 = 32'd9
; 
32'd23851: dataIn1 = 32'd11
; 
32'd23852: dataIn1 = 32'd13
; 
32'd23853: dataIn1 = 32'd15
; 
32'd23854: dataIn1 = 32'd16
; 
32'd23855: dataIn1 = 32'd17
; 
32'd23856: dataIn1 = 32'd18
; 
32'd23857: dataIn1 = 32'd20
; 
32'd23858: dataIn1 = 32'd21
; 
32'd23859: dataIn1 = 32'd25
; 
32'd23860: dataIn1 = 32'd26
; 
32'd23861: dataIn1 = 32'd27
; 
32'd23862: dataIn1 = 32'd31
; 
32'd23863: dataIn1 = 32'd37
; 
32'd23864: dataIn1 = 32'd38
; 
32'd23865: dataIn1 = 32'd39
; 
32'd23866: dataIn1 = 32'd44
; 
32'd23867: dataIn1 = 32'd47
; 
32'd23868: dataIn1 = 32'd53
; 
32'd23869: dataIn1 = 32'd54
; 
32'd23870: dataIn1 = 32'd56
; 
32'd23871: dataIn1 = 32'd57
; 
32'd23872: dataIn1 = 32'd58
; 
32'd23873: dataIn1 = 32'd62
; 
32'd23874: dataIn1 = 32'd63
; 
32'd23875: dataIn1 = 32'd4
; 
32'd23876: dataIn1 = 32'd5
; 
32'd23877: dataIn1 = 32'd6
; 
32'd23878: dataIn1 = 32'd8
; 
32'd23879: dataIn1 = 32'd10
; 
32'd23880: dataIn1 = 32'd11
; 
32'd23881: dataIn1 = 32'd13
; 
32'd23882: dataIn1 = 32'd14
; 
32'd23883: dataIn1 = 32'd17
; 
32'd23884: dataIn1 = 32'd18
; 
32'd23885: dataIn1 = 32'd21
; 
32'd23886: dataIn1 = 32'd28
; 
32'd23887: dataIn1 = 32'd30
; 
32'd23888: dataIn1 = 32'd31
; 
32'd23889: dataIn1 = 32'd33
; 
32'd23890: dataIn1 = 32'd34
; 
32'd23891: dataIn1 = 32'd37
; 
32'd23892: dataIn1 = 32'd43
; 
32'd23893: dataIn1 = 32'd47
; 
32'd23894: dataIn1 = 32'd51
; 
32'd23895: dataIn1 = 32'd53
; 
32'd23896: dataIn1 = 32'd55
; 
32'd23897: dataIn1 = 32'd57
; 
32'd23898: dataIn1 = 32'd58
; 
32'd23899: dataIn1 = 32'd60
; 
32'd23900: dataIn1 = 32'd62
; 
32'd23901: dataIn1 = 32'd0
; 
32'd23902: dataIn1 = 32'd1
; 
32'd23903: dataIn1 = 32'd2
; 
32'd23904: dataIn1 = 32'd3
; 
32'd23905: dataIn1 = 32'd5
; 
32'd23906: dataIn1 = 32'd7
; 
32'd23907: dataIn1 = 32'd11
; 
32'd23908: dataIn1 = 32'd17
; 
32'd23909: dataIn1 = 32'd21
; 
32'd23910: dataIn1 = 32'd22
; 
32'd23911: dataIn1 = 32'd23
; 
32'd23912: dataIn1 = 32'd24
; 
32'd23913: dataIn1 = 32'd27
; 
32'd23914: dataIn1 = 32'd28
; 
32'd23915: dataIn1 = 32'd34
; 
32'd23916: dataIn1 = 32'd37
; 
32'd23917: dataIn1 = 32'd38
; 
32'd23918: dataIn1 = 32'd39
; 
32'd23919: dataIn1 = 32'd40
; 
32'd23920: dataIn1 = 32'd41
; 
32'd23921: dataIn1 = 32'd42
; 
32'd23922: dataIn1 = 32'd43
; 
32'd23923: dataIn1 = 32'd47
; 
32'd23924: dataIn1 = 32'd49
; 
32'd23925: dataIn1 = 32'd50
; 
32'd23926: dataIn1 = 32'd51
; 
32'd23927: dataIn1 = 32'd53
; 
32'd23928: dataIn1 = 32'd54
; 
32'd23929: dataIn1 = 32'd55
; 
32'd23930: dataIn1 = 32'd57
; 
32'd23931: dataIn1 = 32'd58
; 
32'd23932: dataIn1 = 32'd59
; 
32'd23933: dataIn1 = 32'd60
; 
32'd23934: dataIn1 = 32'd61
; 
32'd23935: dataIn1 = 32'd2
; 
32'd23936: dataIn1 = 32'd8
; 
32'd23937: dataIn1 = 32'd9
; 
32'd23938: dataIn1 = 32'd11
; 
32'd23939: dataIn1 = 32'd13
; 
32'd23940: dataIn1 = 32'd14
; 
32'd23941: dataIn1 = 32'd15
; 
32'd23942: dataIn1 = 32'd18
; 
32'd23943: dataIn1 = 32'd22
; 
32'd23944: dataIn1 = 32'd23
; 
32'd23945: dataIn1 = 32'd24
; 
32'd23946: dataIn1 = 32'd25
; 
32'd23947: dataIn1 = 32'd26
; 
32'd23948: dataIn1 = 32'd28
; 
32'd23949: dataIn1 = 32'd30
; 
32'd23950: dataIn1 = 32'd32
; 
32'd23951: dataIn1 = 32'd33
; 
32'd23952: dataIn1 = 32'd35
; 
32'd23953: dataIn1 = 32'd36
; 
32'd23954: dataIn1 = 32'd39
; 
32'd23955: dataIn1 = 32'd41
; 
32'd23956: dataIn1 = 32'd42
; 
32'd23957: dataIn1 = 32'd43
; 
32'd23958: dataIn1 = 32'd46
; 
32'd23959: dataIn1 = 32'd47
; 
32'd23960: dataIn1 = 32'd48
; 
32'd23961: dataIn1 = 32'd52
; 
32'd23962: dataIn1 = 32'd55
; 
32'd23963: dataIn1 = 32'd60
; 
32'd23964: dataIn1 = 32'd0
; 
32'd23965: dataIn1 = 32'd1
; 
32'd23966: dataIn1 = 32'd2
; 
32'd23967: dataIn1 = 32'd3
; 
32'd23968: dataIn1 = 32'd8
; 
32'd23969: dataIn1 = 32'd11
; 
32'd23970: dataIn1 = 32'd13
; 
32'd23971: dataIn1 = 32'd14
; 
32'd23972: dataIn1 = 32'd16
; 
32'd23973: dataIn1 = 32'd17
; 
32'd23974: dataIn1 = 32'd18
; 
32'd23975: dataIn1 = 32'd19
; 
32'd23976: dataIn1 = 32'd21
; 
32'd23977: dataIn1 = 32'd25
; 
32'd23978: dataIn1 = 32'd26
; 
32'd23979: dataIn1 = 32'd29
; 
32'd23980: dataIn1 = 32'd31
; 
32'd23981: dataIn1 = 32'd33
; 
32'd23982: dataIn1 = 32'd34
; 
32'd23983: dataIn1 = 32'd36
; 
32'd23984: dataIn1 = 32'd37
; 
32'd23985: dataIn1 = 32'd40
; 
32'd23986: dataIn1 = 32'd42
; 
32'd23987: dataIn1 = 32'd43
; 
32'd23988: dataIn1 = 32'd44
; 
32'd23989: dataIn1 = 32'd45
; 
32'd23990: dataIn1 = 32'd47
; 
32'd23991: dataIn1 = 32'd49
; 
32'd23992: dataIn1 = 32'd51
; 
32'd23993: dataIn1 = 32'd53
; 
32'd23994: dataIn1 = 32'd55
; 
32'd23995: dataIn1 = 32'd62
; 
32'd23996: dataIn1 = 32'd63
; 
32'd23997: dataIn1 = 32'd0
; 
32'd23998: dataIn1 = 32'd2
; 
32'd23999: dataIn1 = 32'd3
; 
32'd24000: dataIn1 = 32'd4
; 
32'd24001: dataIn1 = 32'd5
; 
32'd24002: dataIn1 = 32'd8
; 
32'd24003: dataIn1 = 32'd17
; 
32'd24004: dataIn1 = 32'd18
; 
32'd24005: dataIn1 = 32'd20
; 
32'd24006: dataIn1 = 32'd23
; 
32'd24007: dataIn1 = 32'd24
; 
32'd24008: dataIn1 = 32'd29
; 
32'd24009: dataIn1 = 32'd33
; 
32'd24010: dataIn1 = 32'd34
; 
32'd24011: dataIn1 = 32'd36
; 
32'd24012: dataIn1 = 32'd37
; 
32'd24013: dataIn1 = 32'd38
; 
32'd24014: dataIn1 = 32'd41
; 
32'd24015: dataIn1 = 32'd43
; 
32'd24016: dataIn1 = 32'd44
; 
32'd24017: dataIn1 = 32'd46
; 
32'd24018: dataIn1 = 32'd48
; 
32'd24019: dataIn1 = 32'd50
; 
32'd24020: dataIn1 = 32'd56
; 
32'd24021: dataIn1 = 32'd60
; 
32'd24022: dataIn1 = 32'd63
; 
32'd24023: dataIn1 = 32'd1
; 
32'd24024: dataIn1 = 32'd4
; 
32'd24025: dataIn1 = 32'd5
; 
32'd24026: dataIn1 = 32'd10
; 
32'd24027: dataIn1 = 32'd11
; 
32'd24028: dataIn1 = 32'd17
; 
32'd24029: dataIn1 = 32'd19
; 
32'd24030: dataIn1 = 32'd20
; 
32'd24031: dataIn1 = 32'd21
; 
32'd24032: dataIn1 = 32'd25
; 
32'd24033: dataIn1 = 32'd26
; 
32'd24034: dataIn1 = 32'd27
; 
32'd24035: dataIn1 = 32'd30
; 
32'd24036: dataIn1 = 32'd32
; 
32'd24037: dataIn1 = 32'd33
; 
32'd24038: dataIn1 = 32'd34
; 
32'd24039: dataIn1 = 32'd35
; 
32'd24040: dataIn1 = 32'd40
; 
32'd24041: dataIn1 = 32'd41
; 
32'd24042: dataIn1 = 32'd43
; 
32'd24043: dataIn1 = 32'd45
; 
32'd24044: dataIn1 = 32'd46
; 
32'd24045: dataIn1 = 32'd51
; 
32'd24046: dataIn1 = 32'd52
; 
32'd24047: dataIn1 = 32'd54
; 
32'd24048: dataIn1 = 32'd57
; 
32'd24049: dataIn1 = 32'd2
; 
32'd24050: dataIn1 = 32'd5
; 
32'd24051: dataIn1 = 32'd7
; 
32'd24052: dataIn1 = 32'd9
; 
32'd24053: dataIn1 = 32'd11
; 
32'd24054: dataIn1 = 32'd13
; 
32'd24055: dataIn1 = 32'd15
; 
32'd24056: dataIn1 = 32'd16
; 
32'd24057: dataIn1 = 32'd17
; 
32'd24058: dataIn1 = 32'd18
; 
32'd24059: dataIn1 = 32'd19
; 
32'd24060: dataIn1 = 32'd21
; 
32'd24061: dataIn1 = 32'd23
; 
32'd24062: dataIn1 = 32'd24
; 
32'd24063: dataIn1 = 32'd25
; 
32'd24064: dataIn1 = 32'd26
; 
32'd24065: dataIn1 = 32'd27
; 
32'd24066: dataIn1 = 32'd31
; 
32'd24067: dataIn1 = 32'd32
; 
32'd24068: dataIn1 = 32'd33
; 
32'd24069: dataIn1 = 32'd34
; 
32'd24070: dataIn1 = 32'd35
; 
32'd24071: dataIn1 = 32'd38
; 
32'd24072: dataIn1 = 32'd40
; 
32'd24073: dataIn1 = 32'd41
; 
32'd24074: dataIn1 = 32'd42
; 
32'd24075: dataIn1 = 32'd44
; 
32'd24076: dataIn1 = 32'd46
; 
32'd24077: dataIn1 = 32'd48
; 
32'd24078: dataIn1 = 32'd49
; 
32'd24079: dataIn1 = 32'd51
; 
32'd24080: dataIn1 = 32'd52
; 
32'd24081: dataIn1 = 32'd54
; 
32'd24082: dataIn1 = 32'd57
; 
32'd24083: dataIn1 = 32'd58
; 
32'd24084: dataIn1 = 32'd59
; 
32'd24085: dataIn1 = 32'd63
; 
32'd24086: dataIn1 = 32'd0
; 
32'd24087: dataIn1 = 32'd1
; 
32'd24088: dataIn1 = 32'd3
; 
32'd24089: dataIn1 = 32'd4
; 
32'd24090: dataIn1 = 32'd9
; 
32'd24091: dataIn1 = 32'd10
; 
32'd24092: dataIn1 = 32'd12
; 
32'd24093: dataIn1 = 32'd14
; 
32'd24094: dataIn1 = 32'd17
; 
32'd24095: dataIn1 = 32'd18
; 
32'd24096: dataIn1 = 32'd19
; 
32'd24097: dataIn1 = 32'd21
; 
32'd24098: dataIn1 = 32'd22
; 
32'd24099: dataIn1 = 32'd23
; 
32'd24100: dataIn1 = 32'd24
; 
32'd24101: dataIn1 = 32'd25
; 
32'd24102: dataIn1 = 32'd27
; 
32'd24103: dataIn1 = 32'd30
; 
32'd24104: dataIn1 = 32'd32
; 
32'd24105: dataIn1 = 32'd36
; 
32'd24106: dataIn1 = 32'd38
; 
32'd24107: dataIn1 = 32'd39
; 
32'd24108: dataIn1 = 32'd42
; 
32'd24109: dataIn1 = 32'd43
; 
32'd24110: dataIn1 = 32'd46
; 
32'd24111: dataIn1 = 32'd47
; 
32'd24112: dataIn1 = 32'd49
; 
32'd24113: dataIn1 = 32'd50
; 
32'd24114: dataIn1 = 32'd51
; 
32'd24115: dataIn1 = 32'd52
; 
32'd24116: dataIn1 = 32'd54
; 
32'd24117: dataIn1 = 32'd57
; 
32'd24118: dataIn1 = 32'd58
; 
32'd24119: dataIn1 = 32'd60
; 
32'd24120: dataIn1 = 32'd61
; 
32'd24121: dataIn1 = 32'd62
; 
32'd24122: dataIn1 = 32'd63
; 
32'd24123: dataIn1 = 32'd2
; 
32'd24124: dataIn1 = 32'd3
; 
32'd24125: dataIn1 = 32'd5
; 
32'd24126: dataIn1 = 32'd6
; 
32'd24127: dataIn1 = 32'd9
; 
32'd24128: dataIn1 = 32'd11
; 
32'd24129: dataIn1 = 32'd13
; 
32'd24130: dataIn1 = 32'd14
; 
32'd24131: dataIn1 = 32'd16
; 
32'd24132: dataIn1 = 32'd17
; 
32'd24133: dataIn1 = 32'd20
; 
32'd24134: dataIn1 = 32'd22
; 
32'd24135: dataIn1 = 32'd23
; 
32'd24136: dataIn1 = 32'd25
; 
32'd24137: dataIn1 = 32'd26
; 
32'd24138: dataIn1 = 32'd27
; 
32'd24139: dataIn1 = 32'd30
; 
32'd24140: dataIn1 = 32'd31
; 
32'd24141: dataIn1 = 32'd33
; 
32'd24142: dataIn1 = 32'd35
; 
32'd24143: dataIn1 = 32'd38
; 
32'd24144: dataIn1 = 32'd42
; 
32'd24145: dataIn1 = 32'd45
; 
32'd24146: dataIn1 = 32'd48
; 
32'd24147: dataIn1 = 32'd54
; 
32'd24148: dataIn1 = 32'd58
; 
32'd24149: dataIn1 = 32'd59
; 
32'd24150: dataIn1 = 32'd61
; 
32'd24151: dataIn1 = 32'd2
; 
32'd24152: dataIn1 = 32'd4
; 
32'd24153: dataIn1 = 32'd6
; 
32'd24154: dataIn1 = 32'd15
; 
32'd24155: dataIn1 = 32'd18
; 
32'd24156: dataIn1 = 32'd22
; 
32'd24157: dataIn1 = 32'd23
; 
32'd24158: dataIn1 = 32'd28
; 
32'd24159: dataIn1 = 32'd29
; 
32'd24160: dataIn1 = 32'd30
; 
32'd24161: dataIn1 = 32'd31
; 
32'd24162: dataIn1 = 32'd38
; 
32'd24163: dataIn1 = 32'd40
; 
32'd24164: dataIn1 = 32'd42
; 
32'd24165: dataIn1 = 32'd43
; 
32'd24166: dataIn1 = 32'd48
; 
32'd24167: dataIn1 = 32'd51
; 
32'd24168: dataIn1 = 32'd52
; 
32'd24169: dataIn1 = 32'd53
; 
32'd24170: dataIn1 = 32'd54
; 
32'd24171: dataIn1 = 32'd56
; 
32'd24172: dataIn1 = 32'd57
; 
32'd24173: dataIn1 = 32'd58
; 
32'd24174: dataIn1 = 32'd60
; 
32'd24175: dataIn1 = 32'd63
; 
32'd24176: dataIn1 = 32'd0
; 
32'd24177: dataIn1 = 32'd4
; 
32'd24178: dataIn1 = 32'd7
; 
32'd24179: dataIn1 = 32'd9
; 
32'd24180: dataIn1 = 32'd12
; 
32'd24181: dataIn1 = 32'd13
; 
32'd24182: dataIn1 = 32'd14
; 
32'd24183: dataIn1 = 32'd15
; 
32'd24184: dataIn1 = 32'd17
; 
32'd24185: dataIn1 = 32'd20
; 
32'd24186: dataIn1 = 32'd24
; 
32'd24187: dataIn1 = 32'd26
; 
32'd24188: dataIn1 = 32'd30
; 
32'd24189: dataIn1 = 32'd32
; 
32'd24190: dataIn1 = 32'd33
; 
32'd24191: dataIn1 = 32'd36
; 
32'd24192: dataIn1 = 32'd37
; 
32'd24193: dataIn1 = 32'd41
; 
32'd24194: dataIn1 = 32'd45
; 
32'd24195: dataIn1 = 32'd46
; 
32'd24196: dataIn1 = 32'd47
; 
32'd24197: dataIn1 = 32'd50
; 
32'd24198: dataIn1 = 32'd51
; 
32'd24199: dataIn1 = 32'd55
; 
32'd24200: dataIn1 = 32'd56
; 
32'd24201: dataIn1 = 32'd57
; 
32'd24202: dataIn1 = 32'd58
; 
32'd24203: dataIn1 = 32'd60
; 
32'd24204: dataIn1 = 32'd62
; 
32'd24205: dataIn1 = 32'd5
; 
32'd24206: dataIn1 = 32'd9
; 
32'd24207: dataIn1 = 32'd11
; 
32'd24208: dataIn1 = 32'd13
; 
32'd24209: dataIn1 = 32'd14
; 
32'd24210: dataIn1 = 32'd17
; 
32'd24211: dataIn1 = 32'd21
; 
32'd24212: dataIn1 = 32'd22
; 
32'd24213: dataIn1 = 32'd23
; 
32'd24214: dataIn1 = 32'd25
; 
32'd24215: dataIn1 = 32'd26
; 
32'd24216: dataIn1 = 32'd29
; 
32'd24217: dataIn1 = 32'd30
; 
32'd24218: dataIn1 = 32'd34
; 
32'd24219: dataIn1 = 32'd35
; 
32'd24220: dataIn1 = 32'd36
; 
32'd24221: dataIn1 = 32'd38
; 
32'd24222: dataIn1 = 32'd40
; 
32'd24223: dataIn1 = 32'd41
; 
32'd24224: dataIn1 = 32'd42
; 
32'd24225: dataIn1 = 32'd45
; 
32'd24226: dataIn1 = 32'd47
; 
32'd24227: dataIn1 = 32'd48
; 
32'd24228: dataIn1 = 32'd49
; 
32'd24229: dataIn1 = 32'd50
; 
32'd24230: dataIn1 = 32'd51
; 
32'd24231: dataIn1 = 32'd57
; 
32'd24232: dataIn1 = 32'd59
; 
32'd24233: dataIn1 = 32'd61
; 
32'd24234: dataIn1 = 32'd62
; 
32'd24235: dataIn1 = 32'd0
; 
32'd24236: dataIn1 = 32'd2
; 
32'd24237: dataIn1 = 32'd4
; 
32'd24238: dataIn1 = 32'd8
; 
32'd24239: dataIn1 = 32'd12
; 
32'd24240: dataIn1 = 32'd13
; 
32'd24241: dataIn1 = 32'd14
; 
32'd24242: dataIn1 = 32'd16
; 
32'd24243: dataIn1 = 32'd18
; 
32'd24244: dataIn1 = 32'd19
; 
32'd24245: dataIn1 = 32'd20
; 
32'd24246: dataIn1 = 32'd21
; 
32'd24247: dataIn1 = 32'd22
; 
32'd24248: dataIn1 = 32'd24
; 
32'd24249: dataIn1 = 32'd27
; 
32'd24250: dataIn1 = 32'd28
; 
32'd24251: dataIn1 = 32'd30
; 
32'd24252: dataIn1 = 32'd31
; 
32'd24253: dataIn1 = 32'd33
; 
32'd24254: dataIn1 = 32'd38
; 
32'd24255: dataIn1 = 32'd40
; 
32'd24256: dataIn1 = 32'd41
; 
32'd24257: dataIn1 = 32'd43
; 
32'd24258: dataIn1 = 32'd45
; 
32'd24259: dataIn1 = 32'd47
; 
32'd24260: dataIn1 = 32'd48
; 
32'd24261: dataIn1 = 32'd49
; 
32'd24262: dataIn1 = 32'd51
; 
32'd24263: dataIn1 = 32'd54
; 
32'd24264: dataIn1 = 32'd61
; 
32'd24265: dataIn1 = 32'd0
; 
32'd24266: dataIn1 = 32'd3
; 
32'd24267: dataIn1 = 32'd5
; 
32'd24268: dataIn1 = 32'd9
; 
32'd24269: dataIn1 = 32'd10
; 
32'd24270: dataIn1 = 32'd11
; 
32'd24271: dataIn1 = 32'd16
; 
32'd24272: dataIn1 = 32'd22
; 
32'd24273: dataIn1 = 32'd23
; 
32'd24274: dataIn1 = 32'd25
; 
32'd24275: dataIn1 = 32'd27
; 
32'd24276: dataIn1 = 32'd28
; 
32'd24277: dataIn1 = 32'd29
; 
32'd24278: dataIn1 = 32'd30
; 
32'd24279: dataIn1 = 32'd31
; 
32'd24280: dataIn1 = 32'd32
; 
32'd24281: dataIn1 = 32'd33
; 
32'd24282: dataIn1 = 32'd35
; 
32'd24283: dataIn1 = 32'd39
; 
32'd24284: dataIn1 = 32'd41
; 
32'd24285: dataIn1 = 32'd43
; 
32'd24286: dataIn1 = 32'd45
; 
32'd24287: dataIn1 = 32'd46
; 
32'd24288: dataIn1 = 32'd48
; 
32'd24289: dataIn1 = 32'd51
; 
32'd24290: dataIn1 = 32'd55
; 
32'd24291: dataIn1 = 32'd56
; 
32'd24292: dataIn1 = 32'd57
; 
32'd24293: dataIn1 = 32'd61
; 
32'd24294: dataIn1 = 32'd62
; 
32'd24295: dataIn1 = 32'd63
; 
32'd24296: dataIn1 = 32'd1
; 
32'd24297: dataIn1 = 32'd5
; 
32'd24298: dataIn1 = 32'd8
; 
32'd24299: dataIn1 = 32'd9
; 
32'd24300: dataIn1 = 32'd11
; 
32'd24301: dataIn1 = 32'd14
; 
32'd24302: dataIn1 = 32'd15
; 
32'd24303: dataIn1 = 32'd17
; 
32'd24304: dataIn1 = 32'd18
; 
32'd24305: dataIn1 = 32'd21
; 
32'd24306: dataIn1 = 32'd26
; 
32'd24307: dataIn1 = 32'd30
; 
32'd24308: dataIn1 = 32'd31
; 
32'd24309: dataIn1 = 32'd34
; 
32'd24310: dataIn1 = 32'd35
; 
32'd24311: dataIn1 = 32'd38
; 
32'd24312: dataIn1 = 32'd40
; 
32'd24313: dataIn1 = 32'd41
; 
32'd24314: dataIn1 = 32'd43
; 
32'd24315: dataIn1 = 32'd45
; 
32'd24316: dataIn1 = 32'd47
; 
32'd24317: dataIn1 = 32'd49
; 
32'd24318: dataIn1 = 32'd50
; 
32'd24319: dataIn1 = 32'd51
; 
32'd24320: dataIn1 = 32'd54
; 
32'd24321: dataIn1 = 32'd55
; 
32'd24322: dataIn1 = 32'd58
; 
32'd24323: dataIn1 = 32'd60
; 
32'd24324: dataIn1 = 32'd0
; 
32'd24325: dataIn1 = 32'd2
; 
32'd24326: dataIn1 = 32'd6
; 
32'd24327: dataIn1 = 32'd7
; 
32'd24328: dataIn1 = 32'd8
; 
32'd24329: dataIn1 = 32'd9
; 
32'd24330: dataIn1 = 32'd11
; 
32'd24331: dataIn1 = 32'd15
; 
32'd24332: dataIn1 = 32'd19
; 
32'd24333: dataIn1 = 32'd21
; 
32'd24334: dataIn1 = 32'd23
; 
32'd24335: dataIn1 = 32'd28
; 
32'd24336: dataIn1 = 32'd29
; 
32'd24337: dataIn1 = 32'd30
; 
32'd24338: dataIn1 = 32'd34
; 
32'd24339: dataIn1 = 32'd35
; 
32'd24340: dataIn1 = 32'd37
; 
32'd24341: dataIn1 = 32'd39
; 
32'd24342: dataIn1 = 32'd40
; 
32'd24343: dataIn1 = 32'd46
; 
32'd24344: dataIn1 = 32'd48
; 
32'd24345: dataIn1 = 32'd49
; 
32'd24346: dataIn1 = 32'd50
; 
32'd24347: dataIn1 = 32'd52
; 
32'd24348: dataIn1 = 32'd53
; 
32'd24349: dataIn1 = 32'd57
; 
32'd24350: dataIn1 = 32'd58
; 
32'd24351: dataIn1 = 32'd59
; 
32'd24352: dataIn1 = 32'd61
; 
32'd24353: dataIn1 = 32'd63
; 
32'd24354: dataIn1 = 32'd1
; 
32'd24355: dataIn1 = 32'd6
; 
32'd24356: dataIn1 = 32'd9
; 
32'd24357: dataIn1 = 32'd12
; 
32'd24358: dataIn1 = 32'd13
; 
32'd24359: dataIn1 = 32'd15
; 
32'd24360: dataIn1 = 32'd16
; 
32'd24361: dataIn1 = 32'd19
; 
32'd24362: dataIn1 = 32'd21
; 
32'd24363: dataIn1 = 32'd23
; 
32'd24364: dataIn1 = 32'd24
; 
32'd24365: dataIn1 = 32'd26
; 
32'd24366: dataIn1 = 32'd28
; 
32'd24367: dataIn1 = 32'd31
; 
32'd24368: dataIn1 = 32'd32
; 
32'd24369: dataIn1 = 32'd34
; 
32'd24370: dataIn1 = 32'd42
; 
32'd24371: dataIn1 = 32'd44
; 
32'd24372: dataIn1 = 32'd45
; 
32'd24373: dataIn1 = 32'd49
; 
32'd24374: dataIn1 = 32'd50
; 
32'd24375: dataIn1 = 32'd53
; 
32'd24376: dataIn1 = 32'd57
; 
32'd24377: dataIn1 = 32'd58
; 
32'd24378: dataIn1 = 32'd59
; 
32'd24379: dataIn1 = 32'd60
; 
32'd24380: dataIn1 = 32'd0
; 
32'd24381: dataIn1 = 32'd1
; 
32'd24382: dataIn1 = 32'd6
; 
32'd24383: dataIn1 = 32'd10
; 
32'd24384: dataIn1 = 32'd18
; 
32'd24385: dataIn1 = 32'd21
; 
32'd24386: dataIn1 = 32'd22
; 
32'd24387: dataIn1 = 32'd23
; 
32'd24388: dataIn1 = 32'd25
; 
32'd24389: dataIn1 = 32'd26
; 
32'd24390: dataIn1 = 32'd34
; 
32'd24391: dataIn1 = 32'd37
; 
32'd24392: dataIn1 = 32'd38
; 
32'd24393: dataIn1 = 32'd39
; 
32'd24394: dataIn1 = 32'd40
; 
32'd24395: dataIn1 = 32'd41
; 
32'd24396: dataIn1 = 32'd44
; 
32'd24397: dataIn1 = 32'd45
; 
32'd24398: dataIn1 = 32'd47
; 
32'd24399: dataIn1 = 32'd48
; 
32'd24400: dataIn1 = 32'd49
; 
32'd24401: dataIn1 = 32'd52
; 
32'd24402: dataIn1 = 32'd57
; 
32'd24403: dataIn1 = 32'd58
; 
32'd24404: dataIn1 = 32'd62
; 
32'd24405: dataIn1 = 32'd63
; 
32'd24406: dataIn1 = 32'd0
; 
32'd24407: dataIn1 = 32'd4
; 
32'd24408: dataIn1 = 32'd5
; 
32'd24409: dataIn1 = 32'd7
; 
32'd24410: dataIn1 = 32'd10
; 
32'd24411: dataIn1 = 32'd14
; 
32'd24412: dataIn1 = 32'd15
; 
32'd24413: dataIn1 = 32'd16
; 
32'd24414: dataIn1 = 32'd18
; 
32'd24415: dataIn1 = 32'd20
; 
32'd24416: dataIn1 = 32'd21
; 
32'd24417: dataIn1 = 32'd25
; 
32'd24418: dataIn1 = 32'd27
; 
32'd24419: dataIn1 = 32'd28
; 
32'd24420: dataIn1 = 32'd29
; 
32'd24421: dataIn1 = 32'd30
; 
32'd24422: dataIn1 = 32'd31
; 
32'd24423: dataIn1 = 32'd35
; 
32'd24424: dataIn1 = 32'd41
; 
32'd24425: dataIn1 = 32'd47
; 
32'd24426: dataIn1 = 32'd52
; 
32'd24427: dataIn1 = 32'd55
; 
32'd24428: dataIn1 = 32'd59
; 
32'd24429: dataIn1 = 32'd60
; 
32'd24430: dataIn1 = 32'd61
; 
32'd24431: dataIn1 = 32'd63
; 
32'd24432: dataIn1 = 32'd0
; 
32'd24433: dataIn1 = 32'd2
; 
32'd24434: dataIn1 = 32'd3
; 
32'd24435: dataIn1 = 32'd6
; 
32'd24436: dataIn1 = 32'd9
; 
32'd24437: dataIn1 = 32'd11
; 
32'd24438: dataIn1 = 32'd12
; 
32'd24439: dataIn1 = 32'd13
; 
32'd24440: dataIn1 = 32'd14
; 
32'd24441: dataIn1 = 32'd15
; 
32'd24442: dataIn1 = 32'd18
; 
32'd24443: dataIn1 = 32'd19
; 
32'd24444: dataIn1 = 32'd23
; 
32'd24445: dataIn1 = 32'd25
; 
32'd24446: dataIn1 = 32'd27
; 
32'd24447: dataIn1 = 32'd28
; 
32'd24448: dataIn1 = 32'd30
; 
32'd24449: dataIn1 = 32'd31
; 
32'd24450: dataIn1 = 32'd33
; 
32'd24451: dataIn1 = 32'd37
; 
32'd24452: dataIn1 = 32'd39
; 
32'd24453: dataIn1 = 32'd41
; 
32'd24454: dataIn1 = 32'd43
; 
32'd24455: dataIn1 = 32'd45
; 
32'd24456: dataIn1 = 32'd46
; 
32'd24457: dataIn1 = 32'd50
; 
32'd24458: dataIn1 = 32'd56
; 
32'd24459: dataIn1 = 32'd58
; 
32'd24460: dataIn1 = 32'd59
; 
32'd24461: dataIn1 = 32'd60
; 
32'd24462: dataIn1 = 32'd61
; 
32'd24463: dataIn1 = 32'd62
; 
32'd24464: dataIn1 = 32'd63
; 
32'd24465: dataIn1 = 32'd2
; 
32'd24466: dataIn1 = 32'd4
; 
32'd24467: dataIn1 = 32'd6
; 
32'd24468: dataIn1 = 32'd7
; 
32'd24469: dataIn1 = 32'd9
; 
32'd24470: dataIn1 = 32'd10
; 
32'd24471: dataIn1 = 32'd11
; 
32'd24472: dataIn1 = 32'd12
; 
32'd24473: dataIn1 = 32'd14
; 
32'd24474: dataIn1 = 32'd17
; 
32'd24475: dataIn1 = 32'd18
; 
32'd24476: dataIn1 = 32'd23
; 
32'd24477: dataIn1 = 32'd25
; 
32'd24478: dataIn1 = 32'd29
; 
32'd24479: dataIn1 = 32'd34
; 
32'd24480: dataIn1 = 32'd35
; 
32'd24481: dataIn1 = 32'd37
; 
32'd24482: dataIn1 = 32'd39
; 
32'd24483: dataIn1 = 32'd40
; 
32'd24484: dataIn1 = 32'd41
; 
32'd24485: dataIn1 = 32'd42
; 
32'd24486: dataIn1 = 32'd43
; 
32'd24487: dataIn1 = 32'd44
; 
32'd24488: dataIn1 = 32'd45
; 
32'd24489: dataIn1 = 32'd47
; 
32'd24490: dataIn1 = 32'd52
; 
32'd24491: dataIn1 = 32'd54
; 
32'd24492: dataIn1 = 32'd55
; 
32'd24493: dataIn1 = 32'd56
; 
32'd24494: dataIn1 = 32'd57
; 
32'd24495: dataIn1 = 32'd60
; 
32'd24496: dataIn1 = 32'd61
; 
32'd24497: dataIn1 = 32'd0
; 
32'd24498: dataIn1 = 32'd1
; 
32'd24499: dataIn1 = 32'd2
; 
32'd24500: dataIn1 = 32'd3
; 
32'd24501: dataIn1 = 32'd5
; 
32'd24502: dataIn1 = 32'd6
; 
32'd24503: dataIn1 = 32'd9
; 
32'd24504: dataIn1 = 32'd11
; 
32'd24505: dataIn1 = 32'd13
; 
32'd24506: dataIn1 = 32'd16
; 
32'd24507: dataIn1 = 32'd18
; 
32'd24508: dataIn1 = 32'd22
; 
32'd24509: dataIn1 = 32'd23
; 
32'd24510: dataIn1 = 32'd24
; 
32'd24511: dataIn1 = 32'd25
; 
32'd24512: dataIn1 = 32'd27
; 
32'd24513: dataIn1 = 32'd29
; 
32'd24514: dataIn1 = 32'd31
; 
32'd24515: dataIn1 = 32'd35
; 
32'd24516: dataIn1 = 32'd39
; 
32'd24517: dataIn1 = 32'd41
; 
32'd24518: dataIn1 = 32'd42
; 
32'd24519: dataIn1 = 32'd43
; 
32'd24520: dataIn1 = 32'd45
; 
32'd24521: dataIn1 = 32'd47
; 
32'd24522: dataIn1 = 32'd48
; 
32'd24523: dataIn1 = 32'd50
; 
32'd24524: dataIn1 = 32'd51
; 
32'd24525: dataIn1 = 32'd54
; 
32'd24526: dataIn1 = 32'd55
; 
32'd24527: dataIn1 = 32'd56
; 
32'd24528: dataIn1 = 32'd57
; 
32'd24529: dataIn1 = 32'd58
; 
32'd24530: dataIn1 = 32'd60
; 
32'd24531: dataIn1 = 32'd61
; 
32'd24532: dataIn1 = 32'd62
; 
32'd24533: dataIn1 = 32'd4
; 
32'd24534: dataIn1 = 32'd5
; 
32'd24535: dataIn1 = 32'd8
; 
32'd24536: dataIn1 = 32'd9
; 
32'd24537: dataIn1 = 32'd13
; 
32'd24538: dataIn1 = 32'd17
; 
32'd24539: dataIn1 = 32'd20
; 
32'd24540: dataIn1 = 32'd23
; 
32'd24541: dataIn1 = 32'd26
; 
32'd24542: dataIn1 = 32'd34
; 
32'd24543: dataIn1 = 32'd35
; 
32'd24544: dataIn1 = 32'd37
; 
32'd24545: dataIn1 = 32'd40
; 
32'd24546: dataIn1 = 32'd41
; 
32'd24547: dataIn1 = 32'd44
; 
32'd24548: dataIn1 = 32'd46
; 
32'd24549: dataIn1 = 32'd50
; 
32'd24550: dataIn1 = 32'd51
; 
32'd24551: dataIn1 = 32'd52
; 
32'd24552: dataIn1 = 32'd53
; 
32'd24553: dataIn1 = 32'd54
; 
32'd24554: dataIn1 = 32'd58
; 
32'd24555: dataIn1 = 32'd59
; 
32'd24556: dataIn1 = 32'd61
; 
32'd24557: dataIn1 = 32'd62
; 
32'd24558: dataIn1 = 32'd63
; 
32'd24559: dataIn1 = 32'd0
; 
32'd24560: dataIn1 = 32'd3
; 
32'd24561: dataIn1 = 32'd5
; 
32'd24562: dataIn1 = 32'd9
; 
32'd24563: dataIn1 = 32'd10
; 
32'd24564: dataIn1 = 32'd11
; 
32'd24565: dataIn1 = 32'd14
; 
32'd24566: dataIn1 = 32'd15
; 
32'd24567: dataIn1 = 32'd16
; 
32'd24568: dataIn1 = 32'd17
; 
32'd24569: dataIn1 = 32'd19
; 
32'd24570: dataIn1 = 32'd26
; 
32'd24571: dataIn1 = 32'd27
; 
32'd24572: dataIn1 = 32'd28
; 
32'd24573: dataIn1 = 32'd30
; 
32'd24574: dataIn1 = 32'd33
; 
32'd24575: dataIn1 = 32'd37
; 
32'd24576: dataIn1 = 32'd39
; 
32'd24577: dataIn1 = 32'd40
; 
32'd24578: dataIn1 = 32'd41
; 
32'd24579: dataIn1 = 32'd44
; 
32'd24580: dataIn1 = 32'd45
; 
32'd24581: dataIn1 = 32'd47
; 
32'd24582: dataIn1 = 32'd48
; 
32'd24583: dataIn1 = 32'd49
; 
32'd24584: dataIn1 = 32'd53
; 
32'd24585: dataIn1 = 32'd54
; 
32'd24586: dataIn1 = 32'd0
; 
32'd24587: dataIn1 = 32'd2
; 
32'd24588: dataIn1 = 32'd3
; 
32'd24589: dataIn1 = 32'd8
; 
32'd24590: dataIn1 = 32'd12
; 
32'd24591: dataIn1 = 32'd14
; 
32'd24592: dataIn1 = 32'd15
; 
32'd24593: dataIn1 = 32'd16
; 
32'd24594: dataIn1 = 32'd17
; 
32'd24595: dataIn1 = 32'd21
; 
32'd24596: dataIn1 = 32'd22
; 
32'd24597: dataIn1 = 32'd23
; 
32'd24598: dataIn1 = 32'd27
; 
32'd24599: dataIn1 = 32'd28
; 
32'd24600: dataIn1 = 32'd31
; 
32'd24601: dataIn1 = 32'd32
; 
32'd24602: dataIn1 = 32'd34
; 
32'd24603: dataIn1 = 32'd35
; 
32'd24604: dataIn1 = 32'd37
; 
32'd24605: dataIn1 = 32'd38
; 
32'd24606: dataIn1 = 32'd41
; 
32'd24607: dataIn1 = 32'd43
; 
32'd24608: dataIn1 = 32'd44
; 
32'd24609: dataIn1 = 32'd46
; 
32'd24610: dataIn1 = 32'd47
; 
32'd24611: dataIn1 = 32'd49
; 
32'd24612: dataIn1 = 32'd50
; 
32'd24613: dataIn1 = 32'd51
; 
32'd24614: dataIn1 = 32'd57
; 
32'd24615: dataIn1 = 32'd60
; 
32'd24616: dataIn1 = 32'd61
; 
32'd24617: dataIn1 = 32'd63
; 
32'd24618: dataIn1 = 32'd1
; 
32'd24619: dataIn1 = 32'd4
; 
32'd24620: dataIn1 = 32'd5
; 
32'd24621: dataIn1 = 32'd6
; 
32'd24622: dataIn1 = 32'd11
; 
32'd24623: dataIn1 = 32'd12
; 
32'd24624: dataIn1 = 32'd13
; 
32'd24625: dataIn1 = 32'd14
; 
32'd24626: dataIn1 = 32'd15
; 
32'd24627: dataIn1 = 32'd16
; 
32'd24628: dataIn1 = 32'd22
; 
32'd24629: dataIn1 = 32'd23
; 
32'd24630: dataIn1 = 32'd24
; 
32'd24631: dataIn1 = 32'd26
; 
32'd24632: dataIn1 = 32'd27
; 
32'd24633: dataIn1 = 32'd28
; 
32'd24634: dataIn1 = 32'd30
; 
32'd24635: dataIn1 = 32'd33
; 
32'd24636: dataIn1 = 32'd36
; 
32'd24637: dataIn1 = 32'd42
; 
32'd24638: dataIn1 = 32'd43
; 
32'd24639: dataIn1 = 32'd44
; 
32'd24640: dataIn1 = 32'd45
; 
32'd24641: dataIn1 = 32'd46
; 
32'd24642: dataIn1 = 32'd47
; 
32'd24643: dataIn1 = 32'd49
; 
32'd24644: dataIn1 = 32'd51
; 
32'd24645: dataIn1 = 32'd54
; 
32'd24646: dataIn1 = 32'd55
; 
32'd24647: dataIn1 = 32'd58
; 
32'd24648: dataIn1 = 32'd59
; 
32'd24649: dataIn1 = 32'd1
; 
32'd24650: dataIn1 = 32'd4
; 
32'd24651: dataIn1 = 32'd7
; 
32'd24652: dataIn1 = 32'd10
; 
32'd24653: dataIn1 = 32'd12
; 
32'd24654: dataIn1 = 32'd13
; 
32'd24655: dataIn1 = 32'd14
; 
32'd24656: dataIn1 = 32'd15
; 
32'd24657: dataIn1 = 32'd16
; 
32'd24658: dataIn1 = 32'd17
; 
32'd24659: dataIn1 = 32'd19
; 
32'd24660: dataIn1 = 32'd25
; 
32'd24661: dataIn1 = 32'd27
; 
32'd24662: dataIn1 = 32'd30
; 
32'd24663: dataIn1 = 32'd32
; 
32'd24664: dataIn1 = 32'd38
; 
32'd24665: dataIn1 = 32'd41
; 
32'd24666: dataIn1 = 32'd43
; 
32'd24667: dataIn1 = 32'd45
; 
32'd24668: dataIn1 = 32'd46
; 
32'd24669: dataIn1 = 32'd47
; 
32'd24670: dataIn1 = 32'd53
; 
32'd24671: dataIn1 = 32'd54
; 
32'd24672: dataIn1 = 32'd55
; 
32'd24673: dataIn1 = 32'd56
; 
32'd24674: dataIn1 = 32'd58
; 
32'd24675: dataIn1 = 32'd59
; 
32'd24676: dataIn1 = 32'd63
; 
32'd24677: dataIn1 = 32'd0
; 
32'd24678: dataIn1 = 32'd1
; 
32'd24679: dataIn1 = 32'd5
; 
32'd24680: dataIn1 = 32'd6
; 
32'd24681: dataIn1 = 32'd8
; 
32'd24682: dataIn1 = 32'd14
; 
32'd24683: dataIn1 = 32'd21
; 
32'd24684: dataIn1 = 32'd23
; 
32'd24685: dataIn1 = 32'd25
; 
32'd24686: dataIn1 = 32'd28
; 
32'd24687: dataIn1 = 32'd29
; 
32'd24688: dataIn1 = 32'd33
; 
32'd24689: dataIn1 = 32'd40
; 
32'd24690: dataIn1 = 32'd41
; 
32'd24691: dataIn1 = 32'd44
; 
32'd24692: dataIn1 = 32'd45
; 
32'd24693: dataIn1 = 32'd50
; 
32'd24694: dataIn1 = 32'd51
; 
32'd24695: dataIn1 = 32'd52
; 
32'd24696: dataIn1 = 32'd56
; 
32'd24697: dataIn1 = 32'd57
; 
32'd24698: dataIn1 = 32'd58
; 
32'd24699: dataIn1 = 32'd59
; 
32'd24700: dataIn1 = 32'd61
; 
32'd24701: dataIn1 = 32'd62
; 
32'd24702: dataIn1 = 32'd63
; 
32'd24703: dataIn1 = 32'd1
; 
32'd24704: dataIn1 = 32'd2
; 
32'd24705: dataIn1 = 32'd3
; 
32'd24706: dataIn1 = 32'd5
; 
32'd24707: dataIn1 = 32'd8
; 
32'd24708: dataIn1 = 32'd10
; 
32'd24709: dataIn1 = 32'd12
; 
32'd24710: dataIn1 = 32'd13
; 
32'd24711: dataIn1 = 32'd14
; 
32'd24712: dataIn1 = 32'd15
; 
32'd24713: dataIn1 = 32'd16
; 
32'd24714: dataIn1 = 32'd18
; 
32'd24715: dataIn1 = 32'd19
; 
32'd24716: dataIn1 = 32'd21
; 
32'd24717: dataIn1 = 32'd23
; 
32'd24718: dataIn1 = 32'd27
; 
32'd24719: dataIn1 = 32'd30
; 
32'd24720: dataIn1 = 32'd32
; 
32'd24721: dataIn1 = 32'd33
; 
32'd24722: dataIn1 = 32'd35
; 
32'd24723: dataIn1 = 32'd36
; 
32'd24724: dataIn1 = 32'd39
; 
32'd24725: dataIn1 = 32'd44
; 
32'd24726: dataIn1 = 32'd46
; 
32'd24727: dataIn1 = 32'd48
; 
32'd24728: dataIn1 = 32'd50
; 
32'd24729: dataIn1 = 32'd51
; 
32'd24730: dataIn1 = 32'd54
; 
32'd24731: dataIn1 = 32'd55
; 
32'd24732: dataIn1 = 32'd56
; 
32'd24733: dataIn1 = 32'd60
; 
32'd24734: dataIn1 = 32'd62
; 
32'd24735: dataIn1 = 32'd3
; 
32'd24736: dataIn1 = 32'd4
; 
32'd24737: dataIn1 = 32'd6
; 
32'd24738: dataIn1 = 32'd8
; 
32'd24739: dataIn1 = 32'd10
; 
32'd24740: dataIn1 = 32'd16
; 
32'd24741: dataIn1 = 32'd19
; 
32'd24742: dataIn1 = 32'd20
; 
32'd24743: dataIn1 = 32'd21
; 
32'd24744: dataIn1 = 32'd24
; 
32'd24745: dataIn1 = 32'd25
; 
32'd24746: dataIn1 = 32'd27
; 
32'd24747: dataIn1 = 32'd30
; 
32'd24748: dataIn1 = 32'd32
; 
32'd24749: dataIn1 = 32'd33
; 
32'd24750: dataIn1 = 32'd36
; 
32'd24751: dataIn1 = 32'd38
; 
32'd24752: dataIn1 = 32'd39
; 
32'd24753: dataIn1 = 32'd40
; 
32'd24754: dataIn1 = 32'd41
; 
32'd24755: dataIn1 = 32'd42
; 
32'd24756: dataIn1 = 32'd44
; 
32'd24757: dataIn1 = 32'd45
; 
32'd24758: dataIn1 = 32'd46
; 
32'd24759: dataIn1 = 32'd50
; 
32'd24760: dataIn1 = 32'd52
; 
32'd24761: dataIn1 = 32'd53
; 
32'd24762: dataIn1 = 32'd55
; 
32'd24763: dataIn1 = 32'd57
; 
32'd24764: dataIn1 = 32'd60
; 
32'd24765: dataIn1 = 32'd61
; 
32'd24766: dataIn1 = 32'd1
; 
32'd24767: dataIn1 = 32'd2
; 
32'd24768: dataIn1 = 32'd3
; 
32'd24769: dataIn1 = 32'd8
; 
32'd24770: dataIn1 = 32'd9
; 
32'd24771: dataIn1 = 32'd10
; 
32'd24772: dataIn1 = 32'd11
; 
32'd24773: dataIn1 = 32'd12
; 
32'd24774: dataIn1 = 32'd13
; 
32'd24775: dataIn1 = 32'd14
; 
32'd24776: dataIn1 = 32'd17
; 
32'd24777: dataIn1 = 32'd20
; 
32'd24778: dataIn1 = 32'd24
; 
32'd24779: dataIn1 = 32'd25
; 
32'd24780: dataIn1 = 32'd28
; 
32'd24781: dataIn1 = 32'd30
; 
32'd24782: dataIn1 = 32'd32
; 
32'd24783: dataIn1 = 32'd33
; 
32'd24784: dataIn1 = 32'd37
; 
32'd24785: dataIn1 = 32'd38
; 
32'd24786: dataIn1 = 32'd45
; 
32'd24787: dataIn1 = 32'd47
; 
32'd24788: dataIn1 = 32'd48
; 
32'd24789: dataIn1 = 32'd55
; 
32'd24790: dataIn1 = 32'd57
; 
32'd24791: dataIn1 = 32'd2
; 
32'd24792: dataIn1 = 32'd3
; 
32'd24793: dataIn1 = 32'd7
; 
32'd24794: dataIn1 = 32'd8
; 
32'd24795: dataIn1 = 32'd9
; 
32'd24796: dataIn1 = 32'd10
; 
32'd24797: dataIn1 = 32'd15
; 
32'd24798: dataIn1 = 32'd18
; 
32'd24799: dataIn1 = 32'd21
; 
32'd24800: dataIn1 = 32'd25
; 
32'd24801: dataIn1 = 32'd28
; 
32'd24802: dataIn1 = 32'd33
; 
32'd24803: dataIn1 = 32'd35
; 
32'd24804: dataIn1 = 32'd36
; 
32'd24805: dataIn1 = 32'd37
; 
32'd24806: dataIn1 = 32'd38
; 
32'd24807: dataIn1 = 32'd39
; 
32'd24808: dataIn1 = 32'd41
; 
32'd24809: dataIn1 = 32'd42
; 
32'd24810: dataIn1 = 32'd43
; 
32'd24811: dataIn1 = 32'd46
; 
32'd24812: dataIn1 = 32'd50
; 
32'd24813: dataIn1 = 32'd54
; 
32'd24814: dataIn1 = 32'd55
; 
32'd24815: dataIn1 = 32'd56
; 
32'd24816: dataIn1 = 32'd57
; 
32'd24817: dataIn1 = 32'd58
; 
32'd24818: dataIn1 = 32'd60
; 
32'd24819: dataIn1 = 32'd61
; 
32'd24820: dataIn1 = 32'd62
; 
32'd24821: dataIn1 = 32'd63
; 
32'd24822: dataIn1 = 32'd0
; 
32'd24823: dataIn1 = 32'd1
; 
32'd24824: dataIn1 = 32'd2
; 
32'd24825: dataIn1 = 32'd5
; 
32'd24826: dataIn1 = 32'd8
; 
32'd24827: dataIn1 = 32'd12
; 
32'd24828: dataIn1 = 32'd14
; 
32'd24829: dataIn1 = 32'd16
; 
32'd24830: dataIn1 = 32'd18
; 
32'd24831: dataIn1 = 32'd22
; 
32'd24832: dataIn1 = 32'd23
; 
32'd24833: dataIn1 = 32'd24
; 
32'd24834: dataIn1 = 32'd26
; 
32'd24835: dataIn1 = 32'd30
; 
32'd24836: dataIn1 = 32'd32
; 
32'd24837: dataIn1 = 32'd35
; 
32'd24838: dataIn1 = 32'd37
; 
32'd24839: dataIn1 = 32'd38
; 
32'd24840: dataIn1 = 32'd39
; 
32'd24841: dataIn1 = 32'd41
; 
32'd24842: dataIn1 = 32'd42
; 
32'd24843: dataIn1 = 32'd43
; 
32'd24844: dataIn1 = 32'd45
; 
32'd24845: dataIn1 = 32'd46
; 
32'd24846: dataIn1 = 32'd47
; 
32'd24847: dataIn1 = 32'd48
; 
32'd24848: dataIn1 = 32'd50
; 
32'd24849: dataIn1 = 32'd54
; 
32'd24850: dataIn1 = 32'd55
; 
32'd24851: dataIn1 = 32'd59
; 
32'd24852: dataIn1 = 32'd60
; 
32'd24853: dataIn1 = 32'd61
; 
32'd24854: dataIn1 = 32'd63
; 
32'd24855: dataIn1 = 32'd1
; 
32'd24856: dataIn1 = 32'd2
; 
32'd24857: dataIn1 = 32'd3
; 
32'd24858: dataIn1 = 32'd7
; 
32'd24859: dataIn1 = 32'd9
; 
32'd24860: dataIn1 = 32'd11
; 
32'd24861: dataIn1 = 32'd12
; 
32'd24862: dataIn1 = 32'd13
; 
32'd24863: dataIn1 = 32'd15
; 
32'd24864: dataIn1 = 32'd16
; 
32'd24865: dataIn1 = 32'd17
; 
32'd24866: dataIn1 = 32'd19
; 
32'd24867: dataIn1 = 32'd25
; 
32'd24868: dataIn1 = 32'd29
; 
32'd24869: dataIn1 = 32'd32
; 
32'd24870: dataIn1 = 32'd34
; 
32'd24871: dataIn1 = 32'd35
; 
32'd24872: dataIn1 = 32'd38
; 
32'd24873: dataIn1 = 32'd45
; 
32'd24874: dataIn1 = 32'd49
; 
32'd24875: dataIn1 = 32'd52
; 
32'd24876: dataIn1 = 32'd54
; 
32'd24877: dataIn1 = 32'd55
; 
32'd24878: dataIn1 = 32'd58
; 
32'd24879: dataIn1 = 32'd61
; 
32'd24880: dataIn1 = 32'd63
; 
32'd24881: dataIn1 = 32'd3
; 
32'd24882: dataIn1 = 32'd7
; 
32'd24883: dataIn1 = 32'd8
; 
32'd24884: dataIn1 = 32'd13
; 
32'd24885: dataIn1 = 32'd15
; 
32'd24886: dataIn1 = 32'd16
; 
32'd24887: dataIn1 = 32'd18
; 
32'd24888: dataIn1 = 32'd19
; 
32'd24889: dataIn1 = 32'd20
; 
32'd24890: dataIn1 = 32'd21
; 
32'd24891: dataIn1 = 32'd24
; 
32'd24892: dataIn1 = 32'd25
; 
32'd24893: dataIn1 = 32'd27
; 
32'd24894: dataIn1 = 32'd29
; 
32'd24895: dataIn1 = 32'd34
; 
32'd24896: dataIn1 = 32'd38
; 
32'd24897: dataIn1 = 32'd39
; 
32'd24898: dataIn1 = 32'd40
; 
32'd24899: dataIn1 = 32'd41
; 
32'd24900: dataIn1 = 32'd43
; 
32'd24901: dataIn1 = 32'd47
; 
32'd24902: dataIn1 = 32'd48
; 
32'd24903: dataIn1 = 32'd49
; 
32'd24904: dataIn1 = 32'd53
; 
32'd24905: dataIn1 = 32'd55
; 
32'd24906: dataIn1 = 32'd59
; 
32'd24907: dataIn1 = 32'd63
; 
32'd24908: dataIn1 = 32'd1
; 
32'd24909: dataIn1 = 32'd3
; 
32'd24910: dataIn1 = 32'd4
; 
32'd24911: dataIn1 = 32'd6
; 
32'd24912: dataIn1 = 32'd8
; 
32'd24913: dataIn1 = 32'd9
; 
32'd24914: dataIn1 = 32'd12
; 
32'd24915: dataIn1 = 32'd14
; 
32'd24916: dataIn1 = 32'd17
; 
32'd24917: dataIn1 = 32'd20
; 
32'd24918: dataIn1 = 32'd25
; 
32'd24919: dataIn1 = 32'd27
; 
32'd24920: dataIn1 = 32'd30
; 
32'd24921: dataIn1 = 32'd31
; 
32'd24922: dataIn1 = 32'd32
; 
32'd24923: dataIn1 = 32'd33
; 
32'd24924: dataIn1 = 32'd34
; 
32'd24925: dataIn1 = 32'd35
; 
32'd24926: dataIn1 = 32'd38
; 
32'd24927: dataIn1 = 32'd41
; 
32'd24928: dataIn1 = 32'd42
; 
32'd24929: dataIn1 = 32'd43
; 
32'd24930: dataIn1 = 32'd44
; 
32'd24931: dataIn1 = 32'd46
; 
32'd24932: dataIn1 = 32'd49
; 
32'd24933: dataIn1 = 32'd52
; 
32'd24934: dataIn1 = 32'd53
; 
32'd24935: dataIn1 = 32'd54
; 
32'd24936: dataIn1 = 32'd55
; 
32'd24937: dataIn1 = 32'd56
; 
32'd24938: dataIn1 = 32'd57
; 
32'd24939: dataIn1 = 32'd58
; 
32'd24940: dataIn1 = 32'd61
; 
32'd24941: dataIn1 = 32'd0
; 
32'd24942: dataIn1 = 32'd1
; 
32'd24943: dataIn1 = 32'd2
; 
32'd24944: dataIn1 = 32'd3
; 
32'd24945: dataIn1 = 32'd4
; 
32'd24946: dataIn1 = 32'd7
; 
32'd24947: dataIn1 = 32'd8
; 
32'd24948: dataIn1 = 32'd12
; 
32'd24949: dataIn1 = 32'd13
; 
32'd24950: dataIn1 = 32'd14
; 
32'd24951: dataIn1 = 32'd17
; 
32'd24952: dataIn1 = 32'd19
; 
32'd24953: dataIn1 = 32'd20
; 
32'd24954: dataIn1 = 32'd23
; 
32'd24955: dataIn1 = 32'd25
; 
32'd24956: dataIn1 = 32'd27
; 
32'd24957: dataIn1 = 32'd28
; 
32'd24958: dataIn1 = 32'd30
; 
32'd24959: dataIn1 = 32'd36
; 
32'd24960: dataIn1 = 32'd37
; 
32'd24961: dataIn1 = 32'd38
; 
32'd24962: dataIn1 = 32'd39
; 
32'd24963: dataIn1 = 32'd41
; 
32'd24964: dataIn1 = 32'd44
; 
32'd24965: dataIn1 = 32'd45
; 
32'd24966: dataIn1 = 32'd47
; 
32'd24967: dataIn1 = 32'd48
; 
32'd24968: dataIn1 = 32'd50
; 
32'd24969: dataIn1 = 32'd51
; 
32'd24970: dataIn1 = 32'd54
; 
32'd24971: dataIn1 = 32'd55
; 
32'd24972: dataIn1 = 32'd56
; 
32'd24973: dataIn1 = 32'd57
; 
32'd24974: dataIn1 = 32'd58
; 
32'd24975: dataIn1 = 32'd60
; 
32'd24976: dataIn1 = 32'd61
; 
32'd24977: dataIn1 = 32'd62
; 
32'd24978: dataIn1 = 32'd0
; 
32'd24979: dataIn1 = 32'd1
; 
32'd24980: dataIn1 = 32'd4
; 
32'd24981: dataIn1 = 32'd6
; 
32'd24982: dataIn1 = 32'd7
; 
32'd24983: dataIn1 = 32'd8
; 
32'd24984: dataIn1 = 32'd9
; 
32'd24985: dataIn1 = 32'd10
; 
32'd24986: dataIn1 = 32'd11
; 
32'd24987: dataIn1 = 32'd12
; 
32'd24988: dataIn1 = 32'd18
; 
32'd24989: dataIn1 = 32'd19
; 
32'd24990: dataIn1 = 32'd23
; 
32'd24991: dataIn1 = 32'd24
; 
32'd24992: dataIn1 = 32'd28
; 
32'd24993: dataIn1 = 32'd30
; 
32'd24994: dataIn1 = 32'd32
; 
32'd24995: dataIn1 = 32'd33
; 
32'd24996: dataIn1 = 32'd35
; 
32'd24997: dataIn1 = 32'd36
; 
32'd24998: dataIn1 = 32'd37
; 
32'd24999: dataIn1 = 32'd39
; 
32'd25000: dataIn1 = 32'd40
; 
32'd25001: dataIn1 = 32'd43
; 
32'd25002: dataIn1 = 32'd45
; 
32'd25003: dataIn1 = 32'd46
; 
32'd25004: dataIn1 = 32'd47
; 
32'd25005: dataIn1 = 32'd48
; 
32'd25006: dataIn1 = 32'd50
; 
32'd25007: dataIn1 = 32'd51
; 
32'd25008: dataIn1 = 32'd53
; 
32'd25009: dataIn1 = 32'd54
; 
32'd25010: dataIn1 = 32'd57
; 
32'd25011: dataIn1 = 32'd61
; 
32'd25012: dataIn1 = 32'd4
; 
32'd25013: dataIn1 = 32'd5
; 
32'd25014: dataIn1 = 32'd6
; 
32'd25015: dataIn1 = 32'd9
; 
32'd25016: dataIn1 = 32'd10
; 
32'd25017: dataIn1 = 32'd11
; 
32'd25018: dataIn1 = 32'd12
; 
32'd25019: dataIn1 = 32'd13
; 
32'd25020: dataIn1 = 32'd18
; 
32'd25021: dataIn1 = 32'd23
; 
32'd25022: dataIn1 = 32'd26
; 
32'd25023: dataIn1 = 32'd27
; 
32'd25024: dataIn1 = 32'd28
; 
32'd25025: dataIn1 = 32'd29
; 
32'd25026: dataIn1 = 32'd30
; 
32'd25027: dataIn1 = 32'd31
; 
32'd25028: dataIn1 = 32'd36
; 
32'd25029: dataIn1 = 32'd39
; 
32'd25030: dataIn1 = 32'd42
; 
32'd25031: dataIn1 = 32'd43
; 
32'd25032: dataIn1 = 32'd44
; 
32'd25033: dataIn1 = 32'd46
; 
32'd25034: dataIn1 = 32'd49
; 
32'd25035: dataIn1 = 32'd50
; 
32'd25036: dataIn1 = 32'd52
; 
32'd25037: dataIn1 = 32'd54
; 
32'd25038: dataIn1 = 32'd55
; 
32'd25039: dataIn1 = 32'd62
; 
32'd25040: dataIn1 = 32'd0
; 
32'd25041: dataIn1 = 32'd1
; 
32'd25042: dataIn1 = 32'd2
; 
32'd25043: dataIn1 = 32'd6
; 
32'd25044: dataIn1 = 32'd7
; 
32'd25045: dataIn1 = 32'd8
; 
32'd25046: dataIn1 = 32'd9
; 
32'd25047: dataIn1 = 32'd10
; 
32'd25048: dataIn1 = 32'd11
; 
32'd25049: dataIn1 = 32'd13
; 
32'd25050: dataIn1 = 32'd14
; 
32'd25051: dataIn1 = 32'd15
; 
32'd25052: dataIn1 = 32'd16
; 
32'd25053: dataIn1 = 32'd21
; 
32'd25054: dataIn1 = 32'd22
; 
32'd25055: dataIn1 = 32'd23
; 
32'd25056: dataIn1 = 32'd25
; 
32'd25057: dataIn1 = 32'd28
; 
32'd25058: dataIn1 = 32'd31
; 
32'd25059: dataIn1 = 32'd34
; 
32'd25060: dataIn1 = 32'd35
; 
32'd25061: dataIn1 = 32'd36
; 
32'd25062: dataIn1 = 32'd37
; 
32'd25063: dataIn1 = 32'd38
; 
32'd25064: dataIn1 = 32'd39
; 
32'd25065: dataIn1 = 32'd40
; 
32'd25066: dataIn1 = 32'd44
; 
32'd25067: dataIn1 = 32'd45
; 
32'd25068: dataIn1 = 32'd46
; 
32'd25069: dataIn1 = 32'd48
; 
32'd25070: dataIn1 = 32'd50
; 
32'd25071: dataIn1 = 32'd51
; 
32'd25072: dataIn1 = 32'd52
; 
32'd25073: dataIn1 = 32'd54
; 
32'd25074: dataIn1 = 32'd56
; 
32'd25075: dataIn1 = 32'd59
; 
32'd25076: dataIn1 = 32'd60
; 
32'd25077: dataIn1 = 32'd0
; 
32'd25078: dataIn1 = 32'd1
; 
32'd25079: dataIn1 = 32'd2
; 
32'd25080: dataIn1 = 32'd3
; 
32'd25081: dataIn1 = 32'd6
; 
32'd25082: dataIn1 = 32'd8
; 
32'd25083: dataIn1 = 32'd10
; 
32'd25084: dataIn1 = 32'd12
; 
32'd25085: dataIn1 = 32'd17
; 
32'd25086: dataIn1 = 32'd19
; 
32'd25087: dataIn1 = 32'd24
; 
32'd25088: dataIn1 = 32'd26
; 
32'd25089: dataIn1 = 32'd27
; 
32'd25090: dataIn1 = 32'd30
; 
32'd25091: dataIn1 = 32'd34
; 
32'd25092: dataIn1 = 32'd35
; 
32'd25093: dataIn1 = 32'd39
; 
32'd25094: dataIn1 = 32'd44
; 
32'd25095: dataIn1 = 32'd45
; 
32'd25096: dataIn1 = 32'd46
; 
32'd25097: dataIn1 = 32'd47
; 
32'd25098: dataIn1 = 32'd48
; 
32'd25099: dataIn1 = 32'd50
; 
32'd25100: dataIn1 = 32'd51
; 
32'd25101: dataIn1 = 32'd52
; 
32'd25102: dataIn1 = 32'd54
; 
32'd25103: dataIn1 = 32'd55
; 
32'd25104: dataIn1 = 32'd56
; 
32'd25105: dataIn1 = 32'd59
; 
32'd25106: dataIn1 = 32'd60
; 
32'd25107: dataIn1 = 32'd61
; 
32'd25108: dataIn1 = 32'd62
; 
32'd25109: dataIn1 = 32'd0
; 
32'd25110: dataIn1 = 32'd2
; 
32'd25111: dataIn1 = 32'd3
; 
32'd25112: dataIn1 = 32'd5
; 
32'd25113: dataIn1 = 32'd7
; 
32'd25114: dataIn1 = 32'd10
; 
32'd25115: dataIn1 = 32'd13
; 
32'd25116: dataIn1 = 32'd26
; 
32'd25117: dataIn1 = 32'd28
; 
32'd25118: dataIn1 = 32'd30
; 
32'd25119: dataIn1 = 32'd31
; 
32'd25120: dataIn1 = 32'd33
; 
32'd25121: dataIn1 = 32'd35
; 
32'd25122: dataIn1 = 32'd37
; 
32'd25123: dataIn1 = 32'd38
; 
32'd25124: dataIn1 = 32'd39
; 
32'd25125: dataIn1 = 32'd40
; 
32'd25126: dataIn1 = 32'd42
; 
32'd25127: dataIn1 = 32'd43
; 
32'd25128: dataIn1 = 32'd46
; 
32'd25129: dataIn1 = 32'd47
; 
32'd25130: dataIn1 = 32'd50
; 
32'd25131: dataIn1 = 32'd51
; 
32'd25132: dataIn1 = 32'd52
; 
32'd25133: dataIn1 = 32'd54
; 
32'd25134: dataIn1 = 32'd55
; 
32'd25135: dataIn1 = 32'd58
; 
32'd25136: dataIn1 = 32'd62
; 
32'd25137: dataIn1 = 32'd63
; 
32'd25138: dataIn1 = 32'd0
; 
32'd25139: dataIn1 = 32'd5
; 
32'd25140: dataIn1 = 32'd6
; 
32'd25141: dataIn1 = 32'd7
; 
32'd25142: dataIn1 = 32'd8
; 
32'd25143: dataIn1 = 32'd9
; 
32'd25144: dataIn1 = 32'd10
; 
32'd25145: dataIn1 = 32'd16
; 
32'd25146: dataIn1 = 32'd17
; 
32'd25147: dataIn1 = 32'd19
; 
32'd25148: dataIn1 = 32'd20
; 
32'd25149: dataIn1 = 32'd22
; 
32'd25150: dataIn1 = 32'd24
; 
32'd25151: dataIn1 = 32'd29
; 
32'd25152: dataIn1 = 32'd30
; 
32'd25153: dataIn1 = 32'd31
; 
32'd25154: dataIn1 = 32'd32
; 
32'd25155: dataIn1 = 32'd33
; 
32'd25156: dataIn1 = 32'd34
; 
32'd25157: dataIn1 = 32'd35
; 
32'd25158: dataIn1 = 32'd37
; 
32'd25159: dataIn1 = 32'd39
; 
32'd25160: dataIn1 = 32'd40
; 
32'd25161: dataIn1 = 32'd41
; 
32'd25162: dataIn1 = 32'd42
; 
32'd25163: dataIn1 = 32'd45
; 
32'd25164: dataIn1 = 32'd46
; 
32'd25165: dataIn1 = 32'd47
; 
32'd25166: dataIn1 = 32'd51
; 
32'd25167: dataIn1 = 32'd52
; 
32'd25168: dataIn1 = 32'd53
; 
32'd25169: dataIn1 = 32'd56
; 
32'd25170: dataIn1 = 32'd59
; 
32'd25171: dataIn1 = 32'd0
; 
32'd25172: dataIn1 = 32'd3
; 
32'd25173: dataIn1 = 32'd4
; 
32'd25174: dataIn1 = 32'd8
; 
32'd25175: dataIn1 = 32'd10
; 
32'd25176: dataIn1 = 32'd12
; 
32'd25177: dataIn1 = 32'd15
; 
32'd25178: dataIn1 = 32'd17
; 
32'd25179: dataIn1 = 32'd18
; 
32'd25180: dataIn1 = 32'd22
; 
32'd25181: dataIn1 = 32'd24
; 
32'd25182: dataIn1 = 32'd25
; 
32'd25183: dataIn1 = 32'd26
; 
32'd25184: dataIn1 = 32'd27
; 
32'd25185: dataIn1 = 32'd29
; 
32'd25186: dataIn1 = 32'd30
; 
32'd25187: dataIn1 = 32'd37
; 
32'd25188: dataIn1 = 32'd39
; 
32'd25189: dataIn1 = 32'd44
; 
32'd25190: dataIn1 = 32'd45
; 
32'd25191: dataIn1 = 32'd48
; 
32'd25192: dataIn1 = 32'd50
; 
32'd25193: dataIn1 = 32'd51
; 
32'd25194: dataIn1 = 32'd52
; 
32'd25195: dataIn1 = 32'd53
; 
32'd25196: dataIn1 = 32'd55
; 
32'd25197: dataIn1 = 32'd57
; 
32'd25198: dataIn1 = 32'd58
; 
32'd25199: dataIn1 = 32'd59
; 
32'd25200: dataIn1 = 32'd60
; 
32'd25201: dataIn1 = 32'd0
; 
32'd25202: dataIn1 = 32'd2
; 
32'd25203: dataIn1 = 32'd4
; 
32'd25204: dataIn1 = 32'd6
; 
32'd25205: dataIn1 = 32'd8
; 
32'd25206: dataIn1 = 32'd10
; 
32'd25207: dataIn1 = 32'd13
; 
32'd25208: dataIn1 = 32'd14
; 
32'd25209: dataIn1 = 32'd16
; 
32'd25210: dataIn1 = 32'd17
; 
32'd25211: dataIn1 = 32'd19
; 
32'd25212: dataIn1 = 32'd24
; 
32'd25213: dataIn1 = 32'd25
; 
32'd25214: dataIn1 = 32'd28
; 
32'd25215: dataIn1 = 32'd29
; 
32'd25216: dataIn1 = 32'd30
; 
32'd25217: dataIn1 = 32'd31
; 
32'd25218: dataIn1 = 32'd32
; 
32'd25219: dataIn1 = 32'd34
; 
32'd25220: dataIn1 = 32'd43
; 
32'd25221: dataIn1 = 32'd44
; 
32'd25222: dataIn1 = 32'd47
; 
32'd25223: dataIn1 = 32'd48
; 
32'd25224: dataIn1 = 32'd49
; 
32'd25225: dataIn1 = 32'd50
; 
32'd25226: dataIn1 = 32'd51
; 
32'd25227: dataIn1 = 32'd53
; 
32'd25228: dataIn1 = 32'd55
; 
32'd25229: dataIn1 = 32'd56
; 
32'd25230: dataIn1 = 32'd57
; 
32'd25231: dataIn1 = 32'd58
; 
32'd25232: dataIn1 = 32'd61
; 
32'd25233: dataIn1 = 32'd1
; 
32'd25234: dataIn1 = 32'd2
; 
32'd25235: dataIn1 = 32'd3
; 
32'd25236: dataIn1 = 32'd6
; 
32'd25237: dataIn1 = 32'd8
; 
32'd25238: dataIn1 = 32'd10
; 
32'd25239: dataIn1 = 32'd15
; 
32'd25240: dataIn1 = 32'd18
; 
32'd25241: dataIn1 = 32'd19
; 
32'd25242: dataIn1 = 32'd24
; 
32'd25243: dataIn1 = 32'd25
; 
32'd25244: dataIn1 = 32'd26
; 
32'd25245: dataIn1 = 32'd27
; 
32'd25246: dataIn1 = 32'd29
; 
32'd25247: dataIn1 = 32'd30
; 
32'd25248: dataIn1 = 32'd31
; 
32'd25249: dataIn1 = 32'd32
; 
32'd25250: dataIn1 = 32'd35
; 
32'd25251: dataIn1 = 32'd39
; 
32'd25252: dataIn1 = 32'd40
; 
32'd25253: dataIn1 = 32'd42
; 
32'd25254: dataIn1 = 32'd43
; 
32'd25255: dataIn1 = 32'd45
; 
32'd25256: dataIn1 = 32'd49
; 
32'd25257: dataIn1 = 32'd50
; 
32'd25258: dataIn1 = 32'd52
; 
32'd25259: dataIn1 = 32'd56
; 
32'd25260: dataIn1 = 32'd59
; 
32'd25261: dataIn1 = 32'd62
; 
32'd25262: dataIn1 = 32'd2
; 
32'd25263: dataIn1 = 32'd4
; 
32'd25264: dataIn1 = 32'd5
; 
32'd25265: dataIn1 = 32'd6
; 
32'd25266: dataIn1 = 32'd10
; 
32'd25267: dataIn1 = 32'd12
; 
32'd25268: dataIn1 = 32'd15
; 
32'd25269: dataIn1 = 32'd17
; 
32'd25270: dataIn1 = 32'd18
; 
32'd25271: dataIn1 = 32'd19
; 
32'd25272: dataIn1 = 32'd24
; 
32'd25273: dataIn1 = 32'd25
; 
32'd25274: dataIn1 = 32'd26
; 
32'd25275: dataIn1 = 32'd33
; 
32'd25276: dataIn1 = 32'd35
; 
32'd25277: dataIn1 = 32'd38
; 
32'd25278: dataIn1 = 32'd40
; 
32'd25279: dataIn1 = 32'd41
; 
32'd25280: dataIn1 = 32'd42
; 
32'd25281: dataIn1 = 32'd44
; 
32'd25282: dataIn1 = 32'd45
; 
32'd25283: dataIn1 = 32'd46
; 
32'd25284: dataIn1 = 32'd49
; 
32'd25285: dataIn1 = 32'd50
; 
32'd25286: dataIn1 = 32'd51
; 
32'd25287: dataIn1 = 32'd53
; 
32'd25288: dataIn1 = 32'd57
; 
32'd25289: dataIn1 = 32'd63
; 
32'd25290: dataIn1 = 32'd0
; 
32'd25291: dataIn1 = 32'd1
; 
32'd25292: dataIn1 = 32'd2
; 
32'd25293: dataIn1 = 32'd3
; 
32'd25294: dataIn1 = 32'd7
; 
32'd25295: dataIn1 = 32'd10
; 
32'd25296: dataIn1 = 32'd11
; 
32'd25297: dataIn1 = 32'd14
; 
32'd25298: dataIn1 = 32'd15
; 
32'd25299: dataIn1 = 32'd16
; 
32'd25300: dataIn1 = 32'd18
; 
32'd25301: dataIn1 = 32'd20
; 
32'd25302: dataIn1 = 32'd23
; 
32'd25303: dataIn1 = 32'd25
; 
32'd25304: dataIn1 = 32'd27
; 
32'd25305: dataIn1 = 32'd28
; 
32'd25306: dataIn1 = 32'd32
; 
32'd25307: dataIn1 = 32'd34
; 
32'd25308: dataIn1 = 32'd35
; 
32'd25309: dataIn1 = 32'd36
; 
32'd25310: dataIn1 = 32'd40
; 
32'd25311: dataIn1 = 32'd41
; 
32'd25312: dataIn1 = 32'd42
; 
32'd25313: dataIn1 = 32'd44
; 
32'd25314: dataIn1 = 32'd47
; 
32'd25315: dataIn1 = 32'd48
; 
32'd25316: dataIn1 = 32'd49
; 
32'd25317: dataIn1 = 32'd50
; 
32'd25318: dataIn1 = 32'd53
; 
32'd25319: dataIn1 = 32'd57
; 
32'd25320: dataIn1 = 32'd59
; 
32'd25321: dataIn1 = 32'd61
; 
32'd25322: dataIn1 = 32'd62
; 
32'd25323: dataIn1 = 32'd0
; 
32'd25324: dataIn1 = 32'd1
; 
32'd25325: dataIn1 = 32'd2
; 
32'd25326: dataIn1 = 32'd5
; 
32'd25327: dataIn1 = 32'd6
; 
32'd25328: dataIn1 = 32'd8
; 
32'd25329: dataIn1 = 32'd10
; 
32'd25330: dataIn1 = 32'd11
; 
32'd25331: dataIn1 = 32'd13
; 
32'd25332: dataIn1 = 32'd17
; 
32'd25333: dataIn1 = 32'd18
; 
32'd25334: dataIn1 = 32'd24
; 
32'd25335: dataIn1 = 32'd25
; 
32'd25336: dataIn1 = 32'd31
; 
32'd25337: dataIn1 = 32'd34
; 
32'd25338: dataIn1 = 32'd35
; 
32'd25339: dataIn1 = 32'd41
; 
32'd25340: dataIn1 = 32'd42
; 
32'd25341: dataIn1 = 32'd43
; 
32'd25342: dataIn1 = 32'd46
; 
32'd25343: dataIn1 = 32'd48
; 
32'd25344: dataIn1 = 32'd50
; 
32'd25345: dataIn1 = 32'd51
; 
32'd25346: dataIn1 = 32'd52
; 
32'd25347: dataIn1 = 32'd55
; 
32'd25348: dataIn1 = 32'd57
; 
32'd25349: dataIn1 = 32'd58
; 
32'd25350: dataIn1 = 32'd60
; 
32'd25351: dataIn1 = 32'd61
; 
32'd25352: dataIn1 = 32'd62
; 
32'd25353: dataIn1 = 32'd63
; 
32'd25354: dataIn1 = 32'd1
; 
32'd25355: dataIn1 = 32'd2
; 
32'd25356: dataIn1 = 32'd4
; 
32'd25357: dataIn1 = 32'd7
; 
32'd25358: dataIn1 = 32'd8
; 
32'd25359: dataIn1 = 32'd11
; 
32'd25360: dataIn1 = 32'd13
; 
32'd25361: dataIn1 = 32'd14
; 
32'd25362: dataIn1 = 32'd15
; 
32'd25363: dataIn1 = 32'd16
; 
32'd25364: dataIn1 = 32'd18
; 
32'd25365: dataIn1 = 32'd21
; 
32'd25366: dataIn1 = 32'd22
; 
32'd25367: dataIn1 = 32'd23
; 
32'd25368: dataIn1 = 32'd25
; 
32'd25369: dataIn1 = 32'd26
; 
32'd25370: dataIn1 = 32'd28
; 
32'd25371: dataIn1 = 32'd29
; 
32'd25372: dataIn1 = 32'd31
; 
32'd25373: dataIn1 = 32'd33
; 
32'd25374: dataIn1 = 32'd35
; 
32'd25375: dataIn1 = 32'd36
; 
32'd25376: dataIn1 = 32'd40
; 
32'd25377: dataIn1 = 32'd42
; 
32'd25378: dataIn1 = 32'd43
; 
32'd25379: dataIn1 = 32'd44
; 
32'd25380: dataIn1 = 32'd49
; 
32'd25381: dataIn1 = 32'd50
; 
32'd25382: dataIn1 = 32'd51
; 
32'd25383: dataIn1 = 32'd52
; 
32'd25384: dataIn1 = 32'd53
; 
32'd25385: dataIn1 = 32'd55
; 
32'd25386: dataIn1 = 32'd56
; 
32'd25387: dataIn1 = 32'd57
; 
32'd25388: dataIn1 = 32'd62
; 
32'd25389: dataIn1 = 32'd0
; 
32'd25390: dataIn1 = 32'd1
; 
32'd25391: dataIn1 = 32'd4
; 
32'd25392: dataIn1 = 32'd5
; 
32'd25393: dataIn1 = 32'd7
; 
32'd25394: dataIn1 = 32'd10
; 
32'd25395: dataIn1 = 32'd11
; 
32'd25396: dataIn1 = 32'd13
; 
32'd25397: dataIn1 = 32'd14
; 
32'd25398: dataIn1 = 32'd18
; 
32'd25399: dataIn1 = 32'd21
; 
32'd25400: dataIn1 = 32'd23
; 
32'd25401: dataIn1 = 32'd26
; 
32'd25402: dataIn1 = 32'd28
; 
32'd25403: dataIn1 = 32'd30
; 
32'd25404: dataIn1 = 32'd33
; 
32'd25405: dataIn1 = 32'd37
; 
32'd25406: dataIn1 = 32'd38
; 
32'd25407: dataIn1 = 32'd39
; 
32'd25408: dataIn1 = 32'd40
; 
32'd25409: dataIn1 = 32'd44
; 
32'd25410: dataIn1 = 32'd45
; 
32'd25411: dataIn1 = 32'd48
; 
32'd25412: dataIn1 = 32'd49
; 
32'd25413: dataIn1 = 32'd53
; 
32'd25414: dataIn1 = 32'd54
; 
32'd25415: dataIn1 = 32'd58
; 
32'd25416: dataIn1 = 32'd60
; 
32'd25417: dataIn1 = 32'd61
; 
32'd25418: dataIn1 = 32'd62
; 
32'd25419: dataIn1 = 32'd63
; 
32'd25420: dataIn1 = 32'd2
; 
32'd25421: dataIn1 = 32'd6
; 
32'd25422: dataIn1 = 32'd8
; 
32'd25423: dataIn1 = 32'd11
; 
32'd25424: dataIn1 = 32'd12
; 
32'd25425: dataIn1 = 32'd13
; 
32'd25426: dataIn1 = 32'd14
; 
32'd25427: dataIn1 = 32'd17
; 
32'd25428: dataIn1 = 32'd18
; 
32'd25429: dataIn1 = 32'd20
; 
32'd25430: dataIn1 = 32'd22
; 
32'd25431: dataIn1 = 32'd23
; 
32'd25432: dataIn1 = 32'd26
; 
32'd25433: dataIn1 = 32'd28
; 
32'd25434: dataIn1 = 32'd30
; 
32'd25435: dataIn1 = 32'd32
; 
32'd25436: dataIn1 = 32'd34
; 
32'd25437: dataIn1 = 32'd35
; 
32'd25438: dataIn1 = 32'd36
; 
32'd25439: dataIn1 = 32'd37
; 
32'd25440: dataIn1 = 32'd38
; 
32'd25441: dataIn1 = 32'd41
; 
32'd25442: dataIn1 = 32'd45
; 
32'd25443: dataIn1 = 32'd46
; 
32'd25444: dataIn1 = 32'd49
; 
32'd25445: dataIn1 = 32'd52
; 
32'd25446: dataIn1 = 32'd53
; 
32'd25447: dataIn1 = 32'd56
; 
32'd25448: dataIn1 = 32'd61
; 
32'd25449: dataIn1 = 32'd62
; 
32'd25450: dataIn1 = 32'd63
; 
32'd25451: dataIn1 = 32'd0
; 
32'd25452: dataIn1 = 32'd1
; 
32'd25453: dataIn1 = 32'd3
; 
32'd25454: dataIn1 = 32'd4
; 
32'd25455: dataIn1 = 32'd6
; 
32'd25456: dataIn1 = 32'd8
; 
32'd25457: dataIn1 = 32'd9
; 
32'd25458: dataIn1 = 32'd10
; 
32'd25459: dataIn1 = 32'd12
; 
32'd25460: dataIn1 = 32'd13
; 
32'd25461: dataIn1 = 32'd16
; 
32'd25462: dataIn1 = 32'd17
; 
32'd25463: dataIn1 = 32'd18
; 
32'd25464: dataIn1 = 32'd19
; 
32'd25465: dataIn1 = 32'd20
; 
32'd25466: dataIn1 = 32'd25
; 
32'd25467: dataIn1 = 32'd29
; 
32'd25468: dataIn1 = 32'd30
; 
32'd25469: dataIn1 = 32'd32
; 
32'd25470: dataIn1 = 32'd34
; 
32'd25471: dataIn1 = 32'd42
; 
32'd25472: dataIn1 = 32'd44
; 
32'd25473: dataIn1 = 32'd45
; 
32'd25474: dataIn1 = 32'd46
; 
32'd25475: dataIn1 = 32'd47
; 
32'd25476: dataIn1 = 32'd48
; 
32'd25477: dataIn1 = 32'd50
; 
32'd25478: dataIn1 = 32'd53
; 
32'd25479: dataIn1 = 32'd54
; 
32'd25480: dataIn1 = 32'd55
; 
32'd25481: dataIn1 = 32'd58
; 
32'd25482: dataIn1 = 32'd59
; 
32'd25483: dataIn1 = 32'd63
; 
32'd25484: dataIn1 = 32'd0
; 
32'd25485: dataIn1 = 32'd1
; 
32'd25486: dataIn1 = 32'd3
; 
32'd25487: dataIn1 = 32'd5
; 
32'd25488: dataIn1 = 32'd6
; 
32'd25489: dataIn1 = 32'd7
; 
32'd25490: dataIn1 = 32'd9
; 
32'd25491: dataIn1 = 32'd13
; 
32'd25492: dataIn1 = 32'd14
; 
32'd25493: dataIn1 = 32'd16
; 
32'd25494: dataIn1 = 32'd17
; 
32'd25495: dataIn1 = 32'd18
; 
32'd25496: dataIn1 = 32'd19
; 
32'd25497: dataIn1 = 32'd20
; 
32'd25498: dataIn1 = 32'd21
; 
32'd25499: dataIn1 = 32'd22
; 
32'd25500: dataIn1 = 32'd25
; 
32'd25501: dataIn1 = 32'd26
; 
32'd25502: dataIn1 = 32'd27
; 
32'd25503: dataIn1 = 32'd29
; 
32'd25504: dataIn1 = 32'd31
; 
32'd25505: dataIn1 = 32'd34
; 
32'd25506: dataIn1 = 32'd37
; 
32'd25507: dataIn1 = 32'd42
; 
32'd25508: dataIn1 = 32'd43
; 
32'd25509: dataIn1 = 32'd45
; 
32'd25510: dataIn1 = 32'd47
; 
32'd25511: dataIn1 = 32'd48
; 
32'd25512: dataIn1 = 32'd50
; 
32'd25513: dataIn1 = 32'd56
; 
32'd25514: dataIn1 = 32'd57
; 
32'd25515: dataIn1 = 32'd59
; 
32'd25516: dataIn1 = 32'd63
; 
32'd25517: dataIn1 = 32'd0
; 
32'd25518: dataIn1 = 32'd3
; 
32'd25519: dataIn1 = 32'd7
; 
32'd25520: dataIn1 = 32'd8
; 
32'd25521: dataIn1 = 32'd11
; 
32'd25522: dataIn1 = 32'd12
; 
32'd25523: dataIn1 = 32'd13
; 
32'd25524: dataIn1 = 32'd17
; 
32'd25525: dataIn1 = 32'd19
; 
32'd25526: dataIn1 = 32'd20
; 
32'd25527: dataIn1 = 32'd23
; 
32'd25528: dataIn1 = 32'd24
; 
32'd25529: dataIn1 = 32'd25
; 
32'd25530: dataIn1 = 32'd28
; 
32'd25531: dataIn1 = 32'd33
; 
32'd25532: dataIn1 = 32'd34
; 
32'd25533: dataIn1 = 32'd35
; 
32'd25534: dataIn1 = 32'd47
; 
32'd25535: dataIn1 = 32'd48
; 
32'd25536: dataIn1 = 32'd49
; 
32'd25537: dataIn1 = 32'd50
; 
32'd25538: dataIn1 = 32'd51
; 
32'd25539: dataIn1 = 32'd52
; 
32'd25540: dataIn1 = 32'd54
; 
32'd25541: dataIn1 = 32'd55
; 
32'd25542: dataIn1 = 32'd56
; 
32'd25543: dataIn1 = 32'd57
; 
32'd25544: dataIn1 = 32'd58
; 
32'd25545: dataIn1 = 32'd60
; 
32'd25546: dataIn1 = 32'd62
; 
32'd25547: dataIn1 = 32'd63
; 
32'd25548: dataIn1 = 32'd3
; 
32'd25549: dataIn1 = 32'd5
; 
32'd25550: dataIn1 = 32'd9
; 
32'd25551: dataIn1 = 32'd10
; 
32'd25552: dataIn1 = 32'd12
; 
32'd25553: dataIn1 = 32'd14
; 
32'd25554: dataIn1 = 32'd17
; 
32'd25555: dataIn1 = 32'd18
; 
32'd25556: dataIn1 = 32'd20
; 
32'd25557: dataIn1 = 32'd22
; 
32'd25558: dataIn1 = 32'd23
; 
32'd25559: dataIn1 = 32'd24
; 
32'd25560: dataIn1 = 32'd26
; 
32'd25561: dataIn1 = 32'd27
; 
32'd25562: dataIn1 = 32'd29
; 
32'd25563: dataIn1 = 32'd30
; 
32'd25564: dataIn1 = 32'd31
; 
32'd25565: dataIn1 = 32'd33
; 
32'd25566: dataIn1 = 32'd34
; 
32'd25567: dataIn1 = 32'd36
; 
32'd25568: dataIn1 = 32'd39
; 
32'd25569: dataIn1 = 32'd40
; 
32'd25570: dataIn1 = 32'd42
; 
32'd25571: dataIn1 = 32'd45
; 
32'd25572: dataIn1 = 32'd46
; 
32'd25573: dataIn1 = 32'd51
; 
32'd25574: dataIn1 = 32'd54
; 
32'd25575: dataIn1 = 32'd55
; 
32'd25576: dataIn1 = 32'd57
; 
32'd25577: dataIn1 = 32'd60
; 
32'd25578: dataIn1 = 32'd61
; 
32'd25579: dataIn1 = 32'd63
; 
32'd25580: dataIn1 = 32'd0
; 
32'd25581: dataIn1 = 32'd3
; 
32'd25582: dataIn1 = 32'd7
; 
32'd25583: dataIn1 = 32'd11
; 
32'd25584: dataIn1 = 32'd12
; 
32'd25585: dataIn1 = 32'd13
; 
32'd25586: dataIn1 = 32'd14
; 
32'd25587: dataIn1 = 32'd16
; 
32'd25588: dataIn1 = 32'd19
; 
32'd25589: dataIn1 = 32'd20
; 
32'd25590: dataIn1 = 32'd25
; 
32'd25591: dataIn1 = 32'd26
; 
32'd25592: dataIn1 = 32'd30
; 
32'd25593: dataIn1 = 32'd34
; 
32'd25594: dataIn1 = 32'd37
; 
32'd25595: dataIn1 = 32'd40
; 
32'd25596: dataIn1 = 32'd42
; 
32'd25597: dataIn1 = 32'd43
; 
32'd25598: dataIn1 = 32'd44
; 
32'd25599: dataIn1 = 32'd46
; 
32'd25600: dataIn1 = 32'd50
; 
32'd25601: dataIn1 = 32'd55
; 
32'd25602: dataIn1 = 32'd57
; 
32'd25603: dataIn1 = 32'd59
; 
32'd25604: dataIn1 = 32'd60
; 
32'd25605: dataIn1 = 32'd61
; 
32'd25606: dataIn1 = 32'd1
; 
32'd25607: dataIn1 = 32'd5
; 
32'd25608: dataIn1 = 32'd6
; 
32'd25609: dataIn1 = 32'd7
; 
32'd25610: dataIn1 = 32'd8
; 
32'd25611: dataIn1 = 32'd10
; 
32'd25612: dataIn1 = 32'd11
; 
32'd25613: dataIn1 = 32'd14
; 
32'd25614: dataIn1 = 32'd15
; 
32'd25615: dataIn1 = 32'd16
; 
32'd25616: dataIn1 = 32'd17
; 
32'd25617: dataIn1 = 32'd18
; 
32'd25618: dataIn1 = 32'd21
; 
32'd25619: dataIn1 = 32'd22
; 
32'd25620: dataIn1 = 32'd23
; 
32'd25621: dataIn1 = 32'd26
; 
32'd25622: dataIn1 = 32'd27
; 
32'd25623: dataIn1 = 32'd28
; 
32'd25624: dataIn1 = 32'd29
; 
32'd25625: dataIn1 = 32'd30
; 
32'd25626: dataIn1 = 32'd31
; 
32'd25627: dataIn1 = 32'd33
; 
32'd25628: dataIn1 = 32'd34
; 
32'd25629: dataIn1 = 32'd36
; 
32'd25630: dataIn1 = 32'd38
; 
32'd25631: dataIn1 = 32'd39
; 
32'd25632: dataIn1 = 32'd41
; 
32'd25633: dataIn1 = 32'd42
; 
32'd25634: dataIn1 = 32'd43
; 
32'd25635: dataIn1 = 32'd44
; 
32'd25636: dataIn1 = 32'd45
; 
32'd25637: dataIn1 = 32'd47
; 
32'd25638: dataIn1 = 32'd49
; 
32'd25639: dataIn1 = 32'd55
; 
32'd25640: dataIn1 = 32'd58
; 
32'd25641: dataIn1 = 32'd59
; 
32'd25642: dataIn1 = 32'd60
; 
32'd25643: dataIn1 = 32'd61
; 
32'd25644: dataIn1 = 32'd63
; 
32'd25645: dataIn1 = 32'd0
; 
32'd25646: dataIn1 = 32'd1
; 
32'd25647: dataIn1 = 32'd2
; 
32'd25648: dataIn1 = 32'd3
; 
32'd25649: dataIn1 = 32'd4
; 
32'd25650: dataIn1 = 32'd7
; 
32'd25651: dataIn1 = 32'd8
; 
32'd25652: dataIn1 = 32'd9
; 
32'd25653: dataIn1 = 32'd17
; 
32'd25654: dataIn1 = 32'd20
; 
32'd25655: dataIn1 = 32'd21
; 
32'd25656: dataIn1 = 32'd22
; 
32'd25657: dataIn1 = 32'd23
; 
32'd25658: dataIn1 = 32'd25
; 
32'd25659: dataIn1 = 32'd26
; 
32'd25660: dataIn1 = 32'd27
; 
32'd25661: dataIn1 = 32'd29
; 
32'd25662: dataIn1 = 32'd30
; 
32'd25663: dataIn1 = 32'd31
; 
32'd25664: dataIn1 = 32'd34
; 
32'd25665: dataIn1 = 32'd35
; 
32'd25666: dataIn1 = 32'd36
; 
32'd25667: dataIn1 = 32'd37
; 
32'd25668: dataIn1 = 32'd38
; 
32'd25669: dataIn1 = 32'd40
; 
32'd25670: dataIn1 = 32'd41
; 
32'd25671: dataIn1 = 32'd42
; 
32'd25672: dataIn1 = 32'd45
; 
32'd25673: dataIn1 = 32'd46
; 
32'd25674: dataIn1 = 32'd48
; 
32'd25675: dataIn1 = 32'd51
; 
32'd25676: dataIn1 = 32'd56
; 
32'd25677: dataIn1 = 32'd57
; 
32'd25678: dataIn1 = 32'd62
; 
32'd25679: dataIn1 = 32'd63
; 
32'd25680: dataIn1 = 32'd0
; 
32'd25681: dataIn1 = 32'd1
; 
32'd25682: dataIn1 = 32'd2
; 
32'd25683: dataIn1 = 32'd5
; 
32'd25684: dataIn1 = 32'd7
; 
32'd25685: dataIn1 = 32'd8
; 
32'd25686: dataIn1 = 32'd10
; 
32'd25687: dataIn1 = 32'd12
; 
32'd25688: dataIn1 = 32'd13
; 
32'd25689: dataIn1 = 32'd14
; 
32'd25690: dataIn1 = 32'd15
; 
32'd25691: dataIn1 = 32'd17
; 
32'd25692: dataIn1 = 32'd18
; 
32'd25693: dataIn1 = 32'd19
; 
32'd25694: dataIn1 = 32'd20
; 
32'd25695: dataIn1 = 32'd22
; 
32'd25696: dataIn1 = 32'd26
; 
32'd25697: dataIn1 = 32'd28
; 
32'd25698: dataIn1 = 32'd29
; 
32'd25699: dataIn1 = 32'd30
; 
32'd25700: dataIn1 = 32'd32
; 
32'd25701: dataIn1 = 32'd35
; 
32'd25702: dataIn1 = 32'd36
; 
32'd25703: dataIn1 = 32'd40
; 
32'd25704: dataIn1 = 32'd41
; 
32'd25705: dataIn1 = 32'd42
; 
32'd25706: dataIn1 = 32'd46
; 
32'd25707: dataIn1 = 32'd48
; 
32'd25708: dataIn1 = 32'd51
; 
32'd25709: dataIn1 = 32'd52
; 
32'd25710: dataIn1 = 32'd54
; 
32'd25711: dataIn1 = 32'd55
; 
32'd25712: dataIn1 = 32'd60
; 
32'd25713: dataIn1 = 32'd61
; 
32'd25714: dataIn1 = 32'd0
; 
32'd25715: dataIn1 = 32'd3
; 
32'd25716: dataIn1 = 32'd4
; 
32'd25717: dataIn1 = 32'd5
; 
32'd25718: dataIn1 = 32'd6
; 
32'd25719: dataIn1 = 32'd10
; 
32'd25720: dataIn1 = 32'd11
; 
32'd25721: dataIn1 = 32'd12
; 
32'd25722: dataIn1 = 32'd16
; 
32'd25723: dataIn1 = 32'd17
; 
32'd25724: dataIn1 = 32'd18
; 
32'd25725: dataIn1 = 32'd20
; 
32'd25726: dataIn1 = 32'd22
; 
32'd25727: dataIn1 = 32'd26
; 
32'd25728: dataIn1 = 32'd27
; 
32'd25729: dataIn1 = 32'd28
; 
32'd25730: dataIn1 = 32'd29
; 
32'd25731: dataIn1 = 32'd31
; 
32'd25732: dataIn1 = 32'd33
; 
32'd25733: dataIn1 = 32'd37
; 
32'd25734: dataIn1 = 32'd40
; 
32'd25735: dataIn1 = 32'd41
; 
32'd25736: dataIn1 = 32'd44
; 
32'd25737: dataIn1 = 32'd50
; 
32'd25738: dataIn1 = 32'd51
; 
32'd25739: dataIn1 = 32'd52
; 
32'd25740: dataIn1 = 32'd54
; 
32'd25741: dataIn1 = 32'd55
; 
32'd25742: dataIn1 = 32'd56
; 
32'd25743: dataIn1 = 32'd57
; 
32'd25744: dataIn1 = 32'd59
; 
32'd25745: dataIn1 = 32'd61
; 
32'd25746: dataIn1 = 32'd62
; 
32'd25747: dataIn1 = 32'd0
; 
32'd25748: dataIn1 = 32'd1
; 
32'd25749: dataIn1 = 32'd2
; 
32'd25750: dataIn1 = 32'd4
; 
32'd25751: dataIn1 = 32'd5
; 
32'd25752: dataIn1 = 32'd8
; 
32'd25753: dataIn1 = 32'd11
; 
32'd25754: dataIn1 = 32'd13
; 
32'd25755: dataIn1 = 32'd18
; 
32'd25756: dataIn1 = 32'd19
; 
32'd25757: dataIn1 = 32'd21
; 
32'd25758: dataIn1 = 32'd22
; 
32'd25759: dataIn1 = 32'd24
; 
32'd25760: dataIn1 = 32'd26
; 
32'd25761: dataIn1 = 32'd27
; 
32'd25762: dataIn1 = 32'd29
; 
32'd25763: dataIn1 = 32'd34
; 
32'd25764: dataIn1 = 32'd35
; 
32'd25765: dataIn1 = 32'd38
; 
32'd25766: dataIn1 = 32'd40
; 
32'd25767: dataIn1 = 32'd42
; 
32'd25768: dataIn1 = 32'd45
; 
32'd25769: dataIn1 = 32'd46
; 
32'd25770: dataIn1 = 32'd48
; 
32'd25771: dataIn1 = 32'd49
; 
32'd25772: dataIn1 = 32'd50
; 
32'd25773: dataIn1 = 32'd52
; 
32'd25774: dataIn1 = 32'd55
; 
32'd25775: dataIn1 = 32'd57
; 
32'd25776: dataIn1 = 32'd59
; 
32'd25777: dataIn1 = 32'd60
; 
32'd25778: dataIn1 = 32'd63
; 
32'd25779: dataIn1 = 32'd3
; 
32'd25780: dataIn1 = 32'd5
; 
32'd25781: dataIn1 = 32'd13
; 
32'd25782: dataIn1 = 32'd17
; 
32'd25783: dataIn1 = 32'd18
; 
32'd25784: dataIn1 = 32'd20
; 
32'd25785: dataIn1 = 32'd21
; 
32'd25786: dataIn1 = 32'd25
; 
32'd25787: dataIn1 = 32'd26
; 
32'd25788: dataIn1 = 32'd27
; 
32'd25789: dataIn1 = 32'd28
; 
32'd25790: dataIn1 = 32'd34
; 
32'd25791: dataIn1 = 32'd36
; 
32'd25792: dataIn1 = 32'd39
; 
32'd25793: dataIn1 = 32'd40
; 
32'd25794: dataIn1 = 32'd42
; 
32'd25795: dataIn1 = 32'd44
; 
32'd25796: dataIn1 = 32'd45
; 
32'd25797: dataIn1 = 32'd47
; 
32'd25798: dataIn1 = 32'd48
; 
32'd25799: dataIn1 = 32'd53
; 
32'd25800: dataIn1 = 32'd54
; 
32'd25801: dataIn1 = 32'd56
; 
32'd25802: dataIn1 = 32'd57
; 
32'd25803: dataIn1 = 32'd59
; 
32'd25804: dataIn1 = 32'd61
; 
32'd25805: dataIn1 = 32'd63
; 
32'd25806: dataIn1 = 32'd; 
32'd25807: dataIn1 = 32'd; 
32'd25808: dataIn1 = 32'd; 
32'd25809: dataIn1 = 32'd; 
32'd25810: dataIn1 = 32'd; 
32'd25811: dataIn1 = 32'd; 
32'd25812: dataIn1 = 32'd; 
32'd25813: dataIn1 = 32'd; 
32'd25814: dataIn1 = 32'd; 
32'd25815: dataIn1 = 32'd; 
32'd25816: dataIn1 = 32'd; 
32'd25817: dataIn1 = 32'd; 
32'd25818: dataIn1 = 32'd; 
32'd25819: dataIn1 = 32'd; 
32'd25820: dataIn1 = 32'd; 
32'd25821: dataIn1 = 32'd; 
32'd25822: dataIn1 = 32'd; 
32'd25823: dataIn1 = 32'd; 
32'd25824: dataIn1 = 32'd; 
32'd25825: dataIn1 = 32'd; 
32'd25826: dataIn1 = 32'd; 
32'd25827: dataIn1 = 32'd; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd77; 
32'd3: dataIn2 = 32'd1; 
32'd4: dataIn2 = 32'd51; 
32'd5: dataIn2 = 32'd78; 
32'd6: dataIn2 = 32'd84; 
32'd7: dataIn2 = 32'd60; 
32'd8: dataIn2 = 32'd94; 
32'd9: dataIn2 = 32'd23; 
32'd10: dataIn2 = 32'd10; 
32'd11: dataIn2 = 32'd22; 
32'd12: dataIn2 = 32'd45; 
32'd13: dataIn2 = 32'd41; 
32'd14: dataIn2 = 32'd94; 
32'd15: dataIn2 = 32'd86; 
32'd16: dataIn2 = 32'd37; 
32'd17: dataIn2 = 32'd60; 
32'd18: dataIn2 = 32'd20; 
32'd19: dataIn2 = 32'd84; 
32'd20: dataIn2 = 32'd41; 
32'd21: dataIn2 = 32'd72; 
32'd22: dataIn2 = 32'd85; 
32'd23: dataIn2 = 32'd80; 
32'd24: dataIn2 = 32'd64; 
32'd25: dataIn2 = 32'd37; 
32'd26: dataIn2 = 32'd1; 
32'd27: dataIn2 = 32'd99; 
32'd28: dataIn2 = 32'd8; 
32'd29: dataIn2 = 32'd87; 
32'd30: dataIn2 = 32'd95; 
32'd31: dataIn2 = 32'd77; 
32'd32: dataIn2 = 32'd88; 
32'd33: dataIn2 = 32'd26; 
32'd34: dataIn2 = 32'd75; 
32'd35: dataIn2 = 32'd70; 
32'd36: dataIn2 = 32'd55; 
32'd37: dataIn2 = 32'd55; 
32'd38: dataIn2 = 32'd53; 
32'd39: dataIn2 = 32'd60; 
32'd40: dataIn2 = 32'd14; 
32'd41: dataIn2 = 32'd87; 
32'd42: dataIn2 = 32'd36; 
32'd43: dataIn2 = 32'd21; 
32'd44: dataIn2 = 32'd66; 
32'd45: dataIn2 = 32'd45; 
32'd46: dataIn2 = 32'd40; 
32'd47: dataIn2 = 32'd61; 
32'd48: dataIn2 = 32'd100; 
32'd49: dataIn2 = 32'd8; 
32'd50: dataIn2 = 32'd60; 
32'd51: dataIn2 = 32'd27; 
32'd52: dataIn2 = 32'd6; 
32'd53: dataIn2 = 32'd70; 
32'd54: dataIn2 = 32'd75; 
32'd55: dataIn2 = 32'd88; 
32'd56: dataIn2 = 32'd26; 
32'd57: dataIn2 = 32'd50; 
32'd58: dataIn2 = 32'd43; 
32'd59: dataIn2 = 32'd84; 
32'd60: dataIn2 = 32'd26; 
32'd61: dataIn2 = 32'd14; 
32'd62: dataIn2 = 32'd78; 
32'd63: dataIn2 = 32'd79; 
32'd64: dataIn2 = 32'd77; 
32'd65: dataIn2 = 32'd78; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd330: dataIn2 = 32'd24; 
32'd331: dataIn2 = 32'd11; 
32'd332: dataIn2 = 32'd91; 
32'd333: dataIn2 = 32'd83; 
32'd334: dataIn2 = 32'd27; 
32'd335: dataIn2 = 32'd95; 
32'd336: dataIn2 = 32'd36; 
32'd337: dataIn2 = 32'd81; 
32'd338: dataIn2 = 32'd23; 
32'd339: dataIn2 = 32'd60; 
32'd340: dataIn2 = 32'd27; 
32'd341: dataIn2 = 32'd64; 
32'd342: dataIn2 = 32'd74; 
32'd343: dataIn2 = 32'd6; 
32'd344: dataIn2 = 32'd58; 
32'd345: dataIn2 = 32'd89; 
32'd346: dataIn2 = 32'd24; 
32'd347: dataIn2 = 32'd58; 
32'd348: dataIn2 = 32'd44; 
32'd349: dataIn2 = 32'd80; 
32'd350: dataIn2 = 32'd10; 
32'd351: dataIn2 = 32'd57; 
32'd352: dataIn2 = 32'd68; 
32'd353: dataIn2 = 32'd83; 
32'd354: dataIn2 = 32'd32; 
32'd355: dataIn2 = 32'd1; 
32'd356: dataIn2 = 32'd58; 
32'd357: dataIn2 = 32'd26; 
32'd358: dataIn2 = 32'd58; 
32'd359: dataIn2 = 32'd64; 
32'd360: dataIn2 = 32'd38; 
32'd361: dataIn2 = 32'd77; 
32'd362: dataIn2 = 32'd31; 
32'd363: dataIn2 = 32'd62; 
32'd364: dataIn2 = 32'd17; 
32'd365: dataIn2 = 32'd58; 
32'd366: dataIn2 = 32'd34; 
32'd367: dataIn2 = 32'd75; 
32'd368: dataIn2 = 32'd14; 
32'd369: dataIn2 = 32'd58; 
32'd370: dataIn2 = 32'd66; 
32'd371: dataIn2 = 32'd30; 
32'd372: dataIn2 = 32'd30; 
32'd373: dataIn2 = 32'd82; 
32'd374: dataIn2 = 32'd7; 
32'd375: dataIn2 = 32'd70; 
32'd376: dataIn2 = 32'd97; 
32'd377: dataIn2 = 32'd76; 
32'd378: dataIn2 = 32'd10; 
32'd379: dataIn2 = 32'd19; 
32'd380: dataIn2 = 32'd100; 
32'd381: dataIn2 = 32'd73; 
32'd382: dataIn2 = 32'd25; 
32'd383: dataIn2 = 32'd85; 
32'd384: dataIn2 = 32'd12; 
32'd385: dataIn2 = 32'd79; 
32'd386: dataIn2 = 32'd19; 
32'd387: dataIn2 = 32'd70; 
32'd388: dataIn2 = 32'd71; 
32'd389: dataIn2 = 32'd92; 
32'd390: dataIn2 = 32'd90; 
32'd391: dataIn2 = 32'd38; 
32'd392: dataIn2 = 32'd24; 
32'd393: dataIn2 = 32'd57; 
32'd394: dataIn2 = 32'd43; 
32'd395: dataIn2 = 32'd24; 
32'd396: dataIn2 = 32'd67; 
32'd397: dataIn2 = 32'd76; 
32'd398: dataIn2 = 32'd12; 
32'd399: dataIn2 = 32'd34; 
32'd400: dataIn2 = 32'd25; 
32'd401: dataIn2 = 32'd78; 
32'd402: dataIn2 = 32'd6; 
32'd403: dataIn2 = 32'd2; 
32'd404: dataIn2 = 32'd28; 
32'd405: dataIn2 = 32'd2; 
32'd406: dataIn2 = 32'd91; 
32'd407: dataIn2 = 32'd3; 
32'd408: dataIn2 = 32'd36; 
32'd409: dataIn2 = 32'd61; 
32'd410: dataIn2 = 32'd45; 
32'd411: dataIn2 = 32'd78; 
32'd412: dataIn2 = 32'd93; 
32'd413: dataIn2 = 32'd28; 
32'd414: dataIn2 = 32'd17; 
32'd415: dataIn2 = 32'd23; 
32'd416: dataIn2 = 32'd93; 
32'd417: dataIn2 = 32'd58; 
32'd418: dataIn2 = 32'd90; 
32'd419: dataIn2 = 32'd37; 
32'd420: dataIn2 = 32'd49; 
32'd421: dataIn2 = 32'd88; 
32'd422: dataIn2 = 32'd94; 
32'd423: dataIn2 = 32'd69; 
32'd424: dataIn2 = 32'd69; 
32'd425: dataIn2 = 32'd69; 
32'd426: dataIn2 = 32'd74; 
32'd427: dataIn2 = 32'd12; 
32'd428: dataIn2 = 32'd69; 
32'd429: dataIn2 = 32'd56; 
32'd430: dataIn2 = 32'd46; 
32'd431: dataIn2 = 32'd56; 
32'd432: dataIn2 = 32'd8; 
32'd433: dataIn2 = 32'd93; 
32'd434: dataIn2 = 32'd86; 
32'd435: dataIn2 = 32'd71; 
32'd436: dataIn2 = 32'd47; 
32'd437: dataIn2 = 32'd29; 
32'd438: dataIn2 = 32'd22; 
32'd439: dataIn2 = 32'd66; 
32'd440: dataIn2 = 32'd2; 
32'd441: dataIn2 = 32'd75; 
32'd442: dataIn2 = 32'd83; 
32'd443: dataIn2 = 32'd39; 
32'd444: dataIn2 = 32'd74; 
32'd445: dataIn2 = 32'd45; 
32'd446: dataIn2 = 32'd22; 
32'd447: dataIn2 = 32'd62; 
32'd448: dataIn2 = 32'd15; 
32'd449: dataIn2 = 32'd43; 
32'd450: dataIn2 = 32'd29; 
32'd451: dataIn2 = 32'd29; 
32'd452: dataIn2 = 32'd9; 
32'd453: dataIn2 = 32'd76; 
32'd454: dataIn2 = 32'd66; 
32'd455: dataIn2 = 32'd40; 
32'd456: dataIn2 = 32'd54; 
32'd457: dataIn2 = 32'd93; 
32'd458: dataIn2 = 32'd13; 
32'd459: dataIn2 = 32'd69; 
32'd460: dataIn2 = 32'd63; 
32'd461: dataIn2 = 32'd69; 
32'd462: dataIn2 = 32'd52; 
32'd463: dataIn2 = 32'd57; 
32'd464: dataIn2 = 32'd60; 
32'd465: dataIn2 = 32'd95; 
32'd466: dataIn2 = 32'd91; 
32'd467: dataIn2 = 32'd74; 
32'd468: dataIn2 = 32'd77; 
32'd469: dataIn2 = 32'd88; 
32'd470: dataIn2 = 32'd13; 
32'd471: dataIn2 = 32'd64; 
32'd472: dataIn2 = 32'd59; 
32'd473: dataIn2 = 32'd86; 
32'd474: dataIn2 = 32'd76; 
32'd475: dataIn2 = 32'd7; 
32'd476: dataIn2 = 32'd28; 
32'd477: dataIn2 = 32'd61; 
32'd478: dataIn2 = 32'd29; 
32'd479: dataIn2 = 32'd26; 
32'd480: dataIn2 = 32'd6; 
32'd481: dataIn2 = 32'd8; 
32'd482: dataIn2 = 32'd43; 
32'd483: dataIn2 = 32'd74; 
32'd484: dataIn2 = 32'd95; 
32'd485: dataIn2 = 32'd49; 
32'd486: dataIn2 = 32'd55; 
32'd487: dataIn2 = 32'd99; 
32'd488: dataIn2 = 32'd79; 
32'd489: dataIn2 = 32'd24; 
32'd490: dataIn2 = 32'd48; 
32'd491: dataIn2 = 32'd19; 
32'd492: dataIn2 = 32'd98; 
32'd493: dataIn2 = 32'd78; 
32'd494: dataIn2 = 32'd7; 
32'd495: dataIn2 = 32'd99; 
32'd496: dataIn2 = 32'd25; 
32'd497: dataIn2 = 32'd14; 
32'd498: dataIn2 = 32'd17; 
32'd499: dataIn2 = 32'd32; 
32'd500: dataIn2 = 32'd58; 
32'd501: dataIn2 = 32'd92; 
32'd502: dataIn2 = 32'd87; 
32'd503: dataIn2 = 32'd77; 
32'd504: dataIn2 = 32'd14; 
32'd505: dataIn2 = 32'd41; 
32'd506: dataIn2 = 32'd77; 
32'd507: dataIn2 = 32'd74; 
32'd508: dataIn2 = 32'd7; 
32'd509: dataIn2 = 32'd29; 
32'd510: dataIn2 = 32'd92; 
32'd511: dataIn2 = 32'd35; 
32'd512: dataIn2 = 32'd14; 
32'd513: dataIn2 = 32'd3; 
32'd514: dataIn2 = 32'd68; 
32'd515: dataIn2 = 32'd13; 
32'd516: dataIn2 = 32'd90; 
32'd517: dataIn2 = 32'd16; 
32'd518: dataIn2 = 32'd82; 
32'd519: dataIn2 = 32'd77; 
32'd520: dataIn2 = 32'd48; 
32'd521: dataIn2 = 32'd29; 
32'd522: dataIn2 = 32'd75; 
32'd523: dataIn2 = 32'd11; 
32'd524: dataIn2 = 32'd9; 
32'd525: dataIn2 = 32'd88; 
32'd526: dataIn2 = 32'd32; 
32'd527: dataIn2 = 32'd88; 
32'd528: dataIn2 = 32'd86; 
32'd529: dataIn2 = 32'd81; 
32'd530: dataIn2 = 32'd21; 
32'd531: dataIn2 = 32'd59; 
32'd532: dataIn2 = 32'd70; 
32'd533: dataIn2 = 32'd52; 
32'd534: dataIn2 = 32'd37; 
32'd535: dataIn2 = 32'd13; 
32'd536: dataIn2 = 32'd8; 
32'd537: dataIn2 = 32'd4; 
32'd538: dataIn2 = 32'd91; 
32'd539: dataIn2 = 32'd77; 
32'd540: dataIn2 = 32'd42; 
32'd541: dataIn2 = 32'd84; 
32'd542: dataIn2 = 32'd67; 
32'd543: dataIn2 = 32'd61; 
32'd544: dataIn2 = 32'd91; 
32'd545: dataIn2 = 32'd10; 
32'd546: dataIn2 = 32'd52; 
32'd547: dataIn2 = 32'd20; 
32'd548: dataIn2 = 32'd50; 
32'd549: dataIn2 = 32'd4; 
32'd550: dataIn2 = 32'd60; 
32'd551: dataIn2 = 32'd22; 
32'd552: dataIn2 = 32'd1; 
32'd553: dataIn2 = 32'd80; 
32'd554: dataIn2 = 32'd69; 
32'd555: dataIn2 = 32'd58; 
32'd556: dataIn2 = 32'd67; 
32'd557: dataIn2 = 32'd31; 
32'd558: dataIn2 = 32'd20; 
32'd559: dataIn2 = 32'd67; 
32'd560: dataIn2 = 32'd34; 
32'd561: dataIn2 = 32'd26; 
32'd562: dataIn2 = 32'd44; 
32'd563: dataIn2 = 32'd0; 
32'd564: dataIn2 = 32'd59; 
32'd565: dataIn2 = 32'd55; 
32'd566: dataIn2 = 32'd43; 
32'd567: dataIn2 = 32'd22; 
32'd568: dataIn2 = 32'd73; 
32'd569: dataIn2 = 32'd72; 
32'd570: dataIn2 = 32'd78; 
32'd571: dataIn2 = 32'd98; 
32'd572: dataIn2 = 32'd74; 
32'd573: dataIn2 = 32'd58; 
32'd574: dataIn2 = 32'd100; 
32'd575: dataIn2 = 32'd65; 
32'd576: dataIn2 = 32'd80; 
32'd577: dataIn2 = 32'd71; 
32'd578: dataIn2 = 32'd60; 
32'd579: dataIn2 = 32'd27; 
32'd580: dataIn2 = 32'd20; 
32'd581: dataIn2 = 32'd40; 
32'd582: dataIn2 = 32'd30; 
32'd583: dataIn2 = 32'd7; 
32'd584: dataIn2 = 32'd83; 
32'd585: dataIn2 = 32'd93; 
32'd586: dataIn2 = 32'd82; 
32'd587: dataIn2 = 32'd38; 
32'd588: dataIn2 = 32'd83; 
32'd589: dataIn2 = 32'd34; 
32'd590: dataIn2 = 32'd100; 
32'd591: dataIn2 = 32'd37; 
32'd592: dataIn2 = 32'd73; 
32'd593: dataIn2 = 32'd20; 
32'd594: dataIn2 = 32'd65; 
32'd595: dataIn2 = 32'd26; 
32'd596: dataIn2 = 32'd86; 
32'd597: dataIn2 = 32'd100; 
32'd598: dataIn2 = 32'd67; 
32'd599: dataIn2 = 32'd23; 
32'd600: dataIn2 = 32'd44; 
32'd601: dataIn2 = 32'd33; 
32'd602: dataIn2 = 32'd62; 
32'd603: dataIn2 = 32'd25; 
32'd604: dataIn2 = 32'd29; 
32'd605: dataIn2 = 32'd18; 
32'd606: dataIn2 = 32'd32; 
32'd607: dataIn2 = 32'd94; 
32'd608: dataIn2 = 32'd24; 
32'd609: dataIn2 = 32'd36; 
32'd610: dataIn2 = 32'd13; 
32'd611: dataIn2 = 32'd33; 
32'd612: dataIn2 = 32'd13; 
32'd613: dataIn2 = 32'd100; 
32'd614: dataIn2 = 32'd65; 
32'd615: dataIn2 = 32'd87; 
32'd616: dataIn2 = 32'd60; 
32'd617: dataIn2 = 32'd24; 
32'd618: dataIn2 = 32'd73; 
32'd619: dataIn2 = 32'd16; 
32'd620: dataIn2 = 32'd8; 
32'd621: dataIn2 = 32'd95; 
32'd622: dataIn2 = 32'd57; 
32'd623: dataIn2 = 32'd0; 
32'd624: dataIn2 = 32'd11; 
32'd625: dataIn2 = 32'd26; 
32'd626: dataIn2 = 32'd73; 
32'd627: dataIn2 = 32'd83; 
32'd628: dataIn2 = 32'd98; 
32'd629: dataIn2 = 32'd23; 
32'd630: dataIn2 = 32'd18; 
32'd631: dataIn2 = 32'd45; 
32'd632: dataIn2 = 32'd55; 
32'd633: dataIn2 = 32'd43; 
32'd634: dataIn2 = 32'd28; 
32'd635: dataIn2 = 32'd59; 
32'd636: dataIn2 = 32'd3; 
32'd637: dataIn2 = 32'd49; 
32'd638: dataIn2 = 32'd17; 
32'd639: dataIn2 = 32'd62; 
32'd640: dataIn2 = 32'd85; 
32'd641: dataIn2 = 32'd37; 
32'd642: dataIn2 = 32'd75; 
32'd643: dataIn2 = 32'd68; 
32'd644: dataIn2 = 32'd52; 
32'd645: dataIn2 = 32'd46; 
32'd646: dataIn2 = 32'd57; 
32'd647: dataIn2 = 32'd56; 
32'd648: dataIn2 = 32'd76; 
32'd649: dataIn2 = 32'd75; 
32'd650: dataIn2 = 32'd7; 
32'd651: dataIn2 = 32'd10; 
32'd652: dataIn2 = 32'd44; 
32'd653: dataIn2 = 32'd38; 
32'd654: dataIn2 = 32'd39; 
32'd655: dataIn2 = 32'd94; 
32'd656: dataIn2 = 32'd42; 
32'd657: dataIn2 = 32'd47; 
32'd658: dataIn2 = 32'd67; 
32'd659: dataIn2 = 32'd77; 
32'd660: dataIn2 = 32'd60; 
32'd661: dataIn2 = 32'd63; 
32'd662: dataIn2 = 32'd15; 
32'd663: dataIn2 = 32'd47; 
32'd664: dataIn2 = 32'd52; 
32'd665: dataIn2 = 32'd56; 
32'd666: dataIn2 = 32'd92; 
32'd667: dataIn2 = 32'd71; 
32'd668: dataIn2 = 32'd83; 
32'd669: dataIn2 = 32'd70; 
32'd670: dataIn2 = 32'd66; 
32'd671: dataIn2 = 32'd57; 
32'd672: dataIn2 = 32'd48; 
32'd673: dataIn2 = 32'd34; 
32'd674: dataIn2 = 32'd57; 
32'd675: dataIn2 = 32'd60; 
32'd676: dataIn2 = 32'd34; 
32'd677: dataIn2 = 32'd75; 
32'd678: dataIn2 = 32'd83; 
32'd679: dataIn2 = 32'd34; 
32'd680: dataIn2 = 32'd100; 
32'd681: dataIn2 = 32'd16; 
32'd682: dataIn2 = 32'd59; 
32'd683: dataIn2 = 32'd55; 
32'd684: dataIn2 = 32'd41; 
32'd685: dataIn2 = 32'd13; 
32'd686: dataIn2 = 32'd98; 
32'd687: dataIn2 = 32'd34; 
32'd688: dataIn2 = 32'd0; 
32'd689: dataIn2 = 32'd44; 
32'd690: dataIn2 = 32'd33; 
32'd691: dataIn2 = 32'd35; 
32'd692: dataIn2 = 32'd37; 
32'd693: dataIn2 = 32'd58; 
32'd694: dataIn2 = 32'd19; 
32'd695: dataIn2 = 32'd67; 
32'd696: dataIn2 = 32'd50; 
32'd697: dataIn2 = 32'd36; 
32'd698: dataIn2 = 32'd18; 
32'd699: dataIn2 = 32'd21; 
32'd700: dataIn2 = 32'd38; 
32'd701: dataIn2 = 32'd48; 
32'd702: dataIn2 = 32'd80; 
32'd703: dataIn2 = 32'd15; 
32'd704: dataIn2 = 32'd35; 
32'd705: dataIn2 = 32'd60; 
32'd706: dataIn2 = 32'd79; 
32'd707: dataIn2 = 32'd48; 
32'd708: dataIn2 = 32'd10; 
32'd709: dataIn2 = 32'd72; 
32'd710: dataIn2 = 32'd54; 
32'd711: dataIn2 = 32'd12; 
32'd712: dataIn2 = 32'd85; 
32'd713: dataIn2 = 32'd43; 
32'd714: dataIn2 = 32'd8; 
32'd715: dataIn2 = 32'd22; 
32'd716: dataIn2 = 32'd1; 
32'd717: dataIn2 = 32'd19; 
32'd718: dataIn2 = 32'd68; 
32'd719: dataIn2 = 32'd70; 
32'd720: dataIn2 = 32'd5; 
32'd721: dataIn2 = 32'd57; 
32'd722: dataIn2 = 32'd69; 
32'd723: dataIn2 = 32'd74; 
32'd724: dataIn2 = 32'd53; 
32'd725: dataIn2 = 32'd55; 
32'd726: dataIn2 = 32'd7; 
32'd727: dataIn2 = 32'd42; 
32'd728: dataIn2 = 32'd63; 
32'd729: dataIn2 = 32'd98; 
32'd730: dataIn2 = 32'd31; 
32'd731: dataIn2 = 32'd94; 
32'd732: dataIn2 = 32'd45; 
32'd733: dataIn2 = 32'd15; 
32'd734: dataIn2 = 32'd60; 
32'd735: dataIn2 = 32'd22; 
32'd736: dataIn2 = 32'd39; 
32'd737: dataIn2 = 32'd45; 
32'd738: dataIn2 = 32'd62; 
32'd739: dataIn2 = 32'd14; 
32'd740: dataIn2 = 32'd91; 
32'd741: dataIn2 = 32'd84; 
32'd742: dataIn2 = 32'd85; 
32'd743: dataIn2 = 32'd31; 
32'd744: dataIn2 = 32'd99; 
32'd745: dataIn2 = 32'd70; 
32'd746: dataIn2 = 32'd15; 
32'd747: dataIn2 = 32'd51; 
32'd748: dataIn2 = 32'd98; 
32'd749: dataIn2 = 32'd96; 
32'd750: dataIn2 = 32'd60; 
32'd751: dataIn2 = 32'd95; 
32'd752: dataIn2 = 32'd66; 
32'd753: dataIn2 = 32'd100; 
32'd754: dataIn2 = 32'd14; 
32'd755: dataIn2 = 32'd89; 
32'd756: dataIn2 = 32'd80; 
32'd757: dataIn2 = 32'd66; 
32'd758: dataIn2 = 32'd7; 
32'd759: dataIn2 = 32'd47; 
32'd760: dataIn2 = 32'd95; 
32'd761: dataIn2 = 32'd7; 
32'd762: dataIn2 = 32'd79; 
32'd763: dataIn2 = 32'd71; 
32'd764: dataIn2 = 32'd56; 
32'd765: dataIn2 = 32'd15; 
32'd766: dataIn2 = 32'd6; 
32'd767: dataIn2 = 32'd12; 
32'd768: dataIn2 = 32'd69; 
32'd769: dataIn2 = 32'd35; 
32'd770: dataIn2 = 32'd26; 
32'd771: dataIn2 = 32'd31; 
32'd772: dataIn2 = 32'd33; 
32'd773: dataIn2 = 32'd69; 
32'd774: dataIn2 = 32'd87; 
32'd775: dataIn2 = 32'd47; 
32'd776: dataIn2 = 32'd100; 
32'd777: dataIn2 = 32'd68; 
32'd778: dataIn2 = 32'd23; 
32'd779: dataIn2 = 32'd38; 
32'd780: dataIn2 = 32'd83; 
32'd781: dataIn2 = 32'd25; 
32'd782: dataIn2 = 32'd81; 
32'd783: dataIn2 = 32'd57; 
32'd784: dataIn2 = 32'd27; 
32'd785: dataIn2 = 32'd99; 
32'd786: dataIn2 = 32'd99; 
32'd787: dataIn2 = 32'd80; 
32'd788: dataIn2 = 32'd58; 
32'd789: dataIn2 = 32'd42; 
32'd790: dataIn2 = 32'd58; 
32'd791: dataIn2 = 32'd98; 
32'd792: dataIn2 = 32'd98; 
32'd793: dataIn2 = 32'd62; 
32'd794: dataIn2 = 32'd30; 
32'd795: dataIn2 = 32'd58; 
32'd796: dataIn2 = 32'd65; 
32'd797: dataIn2 = 32'd63; 
32'd798: dataIn2 = 32'd3; 
32'd799: dataIn2 = 32'd38; 
32'd800: dataIn2 = 32'd88; 
32'd801: dataIn2 = 32'd30; 
32'd802: dataIn2 = 32'd10; 
32'd803: dataIn2 = 32'd100; 
32'd804: dataIn2 = 32'd12; 
32'd805: dataIn2 = 32'd24; 
32'd806: dataIn2 = 32'd83; 
32'd807: dataIn2 = 32'd26; 
32'd808: dataIn2 = 32'd80; 
32'd809: dataIn2 = 32'd78; 
32'd810: dataIn2 = 32'd95; 
32'd811: dataIn2 = 32'd6; 
32'd812: dataIn2 = 32'd78; 
32'd813: dataIn2 = 32'd97; 
32'd814: dataIn2 = 32'd54; 
32'd815: dataIn2 = 32'd51; 
32'd816: dataIn2 = 32'd48; 
32'd817: dataIn2 = 32'd29; 
32'd818: dataIn2 = 32'd31; 
32'd819: dataIn2 = 32'd67; 
32'd820: dataIn2 = 32'd42; 
32'd821: dataIn2 = 32'd5; 
32'd822: dataIn2 = 32'd68; 
32'd823: dataIn2 = 32'd70; 
32'd824: dataIn2 = 32'd9; 
32'd825: dataIn2 = 32'd56; 
32'd826: dataIn2 = 32'd3; 
32'd827: dataIn2 = 32'd45; 
32'd828: dataIn2 = 32'd39; 
32'd829: dataIn2 = 32'd91; 
32'd830: dataIn2 = 32'd43; 
32'd831: dataIn2 = 32'd9; 
32'd832: dataIn2 = 32'd83; 
32'd833: dataIn2 = 32'd33; 
32'd834: dataIn2 = 32'd13; 
32'd835: dataIn2 = 32'd94; 
32'd836: dataIn2 = 32'd12; 
32'd837: dataIn2 = 32'd42; 
32'd838: dataIn2 = 32'd30; 
32'd839: dataIn2 = 32'd79; 
32'd840: dataIn2 = 32'd76; 
32'd841: dataIn2 = 32'd43; 
32'd842: dataIn2 = 32'd7; 
32'd843: dataIn2 = 32'd40; 
32'd844: dataIn2 = 32'd54; 
32'd845: dataIn2 = 32'd97; 
32'd846: dataIn2 = 32'd24; 
32'd847: dataIn2 = 32'd6; 
32'd848: dataIn2 = 32'd37; 
32'd849: dataIn2 = 32'd89; 
32'd850: dataIn2 = 32'd35; 
32'd851: dataIn2 = 32'd65; 
32'd852: dataIn2 = 32'd94; 
32'd853: dataIn2 = 32'd30; 
32'd854: dataIn2 = 32'd24; 
32'd855: dataIn2 = 32'd79; 
32'd856: dataIn2 = 32'd3; 
32'd857: dataIn2 = 32'd86; 
32'd858: dataIn2 = 32'd58; 
32'd859: dataIn2 = 32'd97; 
32'd860: dataIn2 = 32'd4; 
32'd861: dataIn2 = 32'd2; 
32'd862: dataIn2 = 32'd75; 
32'd863: dataIn2 = 32'd6; 
32'd864: dataIn2 = 32'd26; 
32'd865: dataIn2 = 32'd80; 
32'd866: dataIn2 = 32'd46; 
32'd867: dataIn2 = 32'd54; 
32'd868: dataIn2 = 32'd77; 
32'd869: dataIn2 = 32'd95; 
32'd870: dataIn2 = 32'd18; 
32'd871: dataIn2 = 32'd74; 
32'd872: dataIn2 = 32'd19; 
32'd873: dataIn2 = 32'd67; 
32'd874: dataIn2 = 32'd17; 
32'd875: dataIn2 = 32'd67; 
32'd876: dataIn2 = 32'd65; 
32'd877: dataIn2 = 32'd95; 
32'd878: dataIn2 = 32'd3; 
32'd879: dataIn2 = 32'd55; 
32'd880: dataIn2 = 32'd63; 
32'd881: dataIn2 = 32'd68; 
32'd882: dataIn2 = 32'd57; 
32'd883: dataIn2 = 32'd9; 
32'd884: dataIn2 = 32'd21; 
32'd885: dataIn2 = 32'd10; 
32'd886: dataIn2 = 32'd25; 
32'd887: dataIn2 = 32'd52; 
32'd888: dataIn2 = 32'd22; 
32'd889: dataIn2 = 32'd34; 
32'd890: dataIn2 = 32'd37; 
32'd891: dataIn2 = 32'd98; 
32'd892: dataIn2 = 32'd20; 
32'd893: dataIn2 = 32'd22; 
32'd894: dataIn2 = 32'd86; 
32'd895: dataIn2 = 32'd22; 
32'd896: dataIn2 = 32'd64; 
32'd897: dataIn2 = 32'd9; 
32'd898: dataIn2 = 32'd95; 
32'd899: dataIn2 = 32'd69; 
32'd900: dataIn2 = 32'd99; 
32'd901: dataIn2 = 32'd17; 
32'd902: dataIn2 = 32'd14; 
32'd903: dataIn2 = 32'd9; 
32'd904: dataIn2 = 32'd4; 
32'd905: dataIn2 = 32'd0; 
32'd906: dataIn2 = 32'd76; 
32'd907: dataIn2 = 32'd62; 
32'd908: dataIn2 = 32'd87; 
32'd909: dataIn2 = 32'd86; 
32'd910: dataIn2 = 32'd29; 
32'd911: dataIn2 = 32'd43; 
32'd912: dataIn2 = 32'd96; 
32'd913: dataIn2 = 32'd33; 
32'd914: dataIn2 = 32'd100; 
32'd915: dataIn2 = 32'd49; 
32'd916: dataIn2 = 32'd41; 
32'd917: dataIn2 = 32'd40; 
32'd918: dataIn2 = 32'd64; 
32'd919: dataIn2 = 32'd99; 
32'd920: dataIn2 = 32'd40; 
32'd921: dataIn2 = 32'd30; 
32'd922: dataIn2 = 32'd17; 
32'd923: dataIn2 = 32'd28; 
32'd924: dataIn2 = 32'd13; 
32'd925: dataIn2 = 32'd30; 
32'd926: dataIn2 = 32'd55; 
32'd927: dataIn2 = 32'd81; 
32'd928: dataIn2 = 32'd41; 
32'd929: dataIn2 = 32'd56; 
32'd930: dataIn2 = 32'd36; 
32'd931: dataIn2 = 32'd92; 
32'd932: dataIn2 = 32'd35; 
32'd933: dataIn2 = 32'd72; 
32'd934: dataIn2 = 32'd32; 
32'd935: dataIn2 = 32'd47; 
32'd936: dataIn2 = 32'd75; 
32'd937: dataIn2 = 32'd4; 
32'd938: dataIn2 = 32'd28; 
32'd939: dataIn2 = 32'd19; 
32'd940: dataIn2 = 32'd3; 
32'd941: dataIn2 = 32'd25; 
32'd942: dataIn2 = 32'd54; 
32'd943: dataIn2 = 32'd44; 
32'd944: dataIn2 = 32'd22; 
32'd945: dataIn2 = 32'd86; 
32'd946: dataIn2 = 32'd41; 
32'd947: dataIn2 = 32'd28; 
32'd948: dataIn2 = 32'd92; 
32'd949: dataIn2 = 32'd35; 
32'd950: dataIn2 = 32'd100; 
32'd951: dataIn2 = 32'd28; 
32'd952: dataIn2 = 32'd12; 
32'd953: dataIn2 = 32'd74; 
32'd954: dataIn2 = 32'd57; 
32'd955: dataIn2 = 32'd1; 
32'd956: dataIn2 = 32'd66; 
32'd957: dataIn2 = 32'd88; 
32'd958: dataIn2 = 32'd94; 
32'd959: dataIn2 = 32'd92; 
32'd960: dataIn2 = 32'd69; 
32'd961: dataIn2 = 32'd79; 
32'd962: dataIn2 = 32'd35; 
32'd963: dataIn2 = 32'd42; 
32'd964: dataIn2 = 32'd89; 
32'd965: dataIn2 = 32'd69; 
32'd966: dataIn2 = 32'd93; 
32'd967: dataIn2 = 32'd26; 
32'd968: dataIn2 = 32'd84; 
32'd969: dataIn2 = 32'd49; 
32'd970: dataIn2 = 32'd65; 
32'd971: dataIn2 = 32'd100; 
32'd972: dataIn2 = 32'd54; 
32'd973: dataIn2 = 32'd77; 
32'd974: dataIn2 = 32'd32; 
32'd975: dataIn2 = 32'd53; 
32'd976: dataIn2 = 32'd96; 
32'd977: dataIn2 = 32'd62; 
32'd978: dataIn2 = 32'd72; 
32'd979: dataIn2 = 32'd30; 
32'd980: dataIn2 = 32'd70; 
32'd981: dataIn2 = 32'd80; 
32'd982: dataIn2 = 32'd6; 
32'd983: dataIn2 = 32'd2; 
32'd984: dataIn2 = 32'd55; 
32'd985: dataIn2 = 32'd79; 
32'd986: dataIn2 = 32'd96; 
32'd987: dataIn2 = 32'd61; 
32'd988: dataIn2 = 32'd5; 
32'd989: dataIn2 = 32'd79; 
32'd990: dataIn2 = 32'd34; 
32'd991: dataIn2 = 32'd96; 
32'd992: dataIn2 = 32'd81; 
32'd993: dataIn2 = 32'd100; 
32'd994: dataIn2 = 32'd73; 
32'd995: dataIn2 = 32'd50; 
32'd996: dataIn2 = 32'd63; 
32'd997: dataIn2 = 32'd80; 
32'd998: dataIn2 = 32'd27; 
32'd999: dataIn2 = 32'd40; 
32'd1000: dataIn2 = 32'd24; 
32'd1001: dataIn2 = 32'd48; 
32'd1002: dataIn2 = 32'd71; 
32'd1003: dataIn2 = 32'd24; 
32'd1004: dataIn2 = 32'd72; 
32'd1005: dataIn2 = 32'd42; 
32'd1006: dataIn2 = 32'd64; 
32'd1007: dataIn2 = 32'd99; 
32'd1008: dataIn2 = 32'd64; 
32'd1009: dataIn2 = 32'd49; 
32'd1010: dataIn2 = 32'd67; 
32'd1011: dataIn2 = 32'd60; 
32'd1012: dataIn2 = 32'd14; 
32'd1013: dataIn2 = 32'd10; 
32'd1014: dataIn2 = 32'd53; 
32'd1015: dataIn2 = 32'd62; 
32'd1016: dataIn2 = 32'd81; 
32'd1017: dataIn2 = 32'd73; 
32'd1018: dataIn2 = 32'd13; 
32'd1019: dataIn2 = 32'd92; 
32'd1020: dataIn2 = 32'd73; 
32'd1021: dataIn2 = 32'd62; 
32'd1022: dataIn2 = 32'd36; 
32'd1023: dataIn2 = 32'd88; 
32'd1024: dataIn2 = 32'd100; 
32'd1025: dataIn2 = 32'd5; 
32'd1026: dataIn2 = 32'd27; 
32'd1027: dataIn2 = 32'd85; 
32'd1028: dataIn2 = 32'd96; 
32'd1029: dataIn2 = 32'd9; 
32'd1030: dataIn2 = 32'd47; 
32'd1031: dataIn2 = 32'd3; 
32'd1032: dataIn2 = 32'd12; 
32'd1033: dataIn2 = 32'd29; 
32'd1034: dataIn2 = 32'd96; 
32'd1035: dataIn2 = 32'd76; 
32'd1036: dataIn2 = 32'd75; 
32'd1037: dataIn2 = 32'd83; 
32'd1038: dataIn2 = 32'd73; 
32'd1039: dataIn2 = 32'd83; 
32'd1040: dataIn2 = 32'd44; 
32'd1041: dataIn2 = 32'd57; 
32'd1042: dataIn2 = 32'd83; 
32'd1043: dataIn2 = 32'd25; 
32'd1044: dataIn2 = 32'd5; 
32'd1045: dataIn2 = 32'd43; 
32'd1046: dataIn2 = 32'd7; 
32'd1047: dataIn2 = 32'd10; 
32'd1048: dataIn2 = 32'd46; 
32'd1049: dataIn2 = 32'd6; 
32'd1050: dataIn2 = 32'd41; 
32'd1051: dataIn2 = 32'd2; 
32'd1052: dataIn2 = 32'd88; 
32'd1053: dataIn2 = 32'd57; 
32'd1054: dataIn2 = 32'd26; 
32'd1055: dataIn2 = 32'd42; 
32'd1056: dataIn2 = 32'd44; 
32'd1057: dataIn2 = 32'd90; 
32'd1058: dataIn2 = 32'd7; 
32'd1059: dataIn2 = 32'd72; 
32'd1060: dataIn2 = 32'd37; 
32'd1061: dataIn2 = 32'd24; 
32'd1062: dataIn2 = 32'd22; 
32'd1063: dataIn2 = 32'd68; 
32'd1064: dataIn2 = 32'd77; 
32'd1065: dataIn2 = 32'd54; 
32'd1066: dataIn2 = 32'd48; 
32'd1067: dataIn2 = 32'd71; 
32'd1068: dataIn2 = 32'd75; 
32'd1069: dataIn2 = 32'd53; 
32'd1070: dataIn2 = 32'd3; 
32'd1071: dataIn2 = 32'd89; 
32'd1072: dataIn2 = 32'd13; 
32'd1073: dataIn2 = 32'd67; 
32'd1074: dataIn2 = 32'd77; 
32'd1075: dataIn2 = 32'd23; 
32'd1076: dataIn2 = 32'd12; 
32'd1077: dataIn2 = 32'd13; 
32'd1078: dataIn2 = 32'd12; 
32'd1079: dataIn2 = 32'd68; 
32'd1080: dataIn2 = 32'd74; 
32'd1081: dataIn2 = 32'd43; 
32'd1082: dataIn2 = 32'd87; 
32'd1083: dataIn2 = 32'd80; 
32'd1084: dataIn2 = 32'd28; 
32'd1085: dataIn2 = 32'd11; 
32'd1086: dataIn2 = 32'd61; 
32'd1087: dataIn2 = 32'd93; 
32'd1088: dataIn2 = 32'd92; 
32'd1089: dataIn2 = 32'd4; 
32'd1090: dataIn2 = 32'd2; 
32'd1091: dataIn2 = 32'd16; 
32'd1092: dataIn2 = 32'd51; 
32'd1093: dataIn2 = 32'd10; 
32'd1094: dataIn2 = 32'd21; 
32'd1095: dataIn2 = 32'd28; 
32'd1096: dataIn2 = 32'd6; 
32'd1097: dataIn2 = 32'd1; 
32'd1098: dataIn2 = 32'd39; 
32'd1099: dataIn2 = 32'd70; 
32'd1100: dataIn2 = 32'd66; 
32'd1101: dataIn2 = 32'd6; 
32'd1102: dataIn2 = 32'd87; 
32'd1103: dataIn2 = 32'd0; 
32'd1104: dataIn2 = 32'd38; 
32'd1105: dataIn2 = 32'd61; 
32'd1106: dataIn2 = 32'd69; 
32'd1107: dataIn2 = 32'd35; 
32'd1108: dataIn2 = 32'd21; 
32'd1109: dataIn2 = 32'd97; 
32'd1110: dataIn2 = 32'd66; 
32'd1111: dataIn2 = 32'd2; 
32'd1112: dataIn2 = 32'd69; 
32'd1113: dataIn2 = 32'd7; 
32'd1114: dataIn2 = 32'd32; 
32'd1115: dataIn2 = 32'd58; 
32'd1116: dataIn2 = 32'd52; 
32'd1117: dataIn2 = 32'd70; 
32'd1118: dataIn2 = 32'd8; 
32'd1119: dataIn2 = 32'd87; 
32'd1120: dataIn2 = 32'd25; 
32'd1121: dataIn2 = 32'd7; 
32'd1122: dataIn2 = 32'd20; 
32'd1123: dataIn2 = 32'd4; 
32'd1124: dataIn2 = 32'd59; 
32'd1125: dataIn2 = 32'd89; 
32'd1126: dataIn2 = 32'd24; 
32'd1127: dataIn2 = 32'd50; 
32'd1128: dataIn2 = 32'd72; 
32'd1129: dataIn2 = 32'd40; 
32'd1130: dataIn2 = 32'd46; 
32'd1131: dataIn2 = 32'd87; 
32'd1132: dataIn2 = 32'd61; 
32'd1133: dataIn2 = 32'd54; 
32'd1134: dataIn2 = 32'd5; 
32'd1135: dataIn2 = 32'd28; 
32'd1136: dataIn2 = 32'd5; 
32'd1137: dataIn2 = 32'd27; 
32'd1138: dataIn2 = 32'd93; 
32'd1139: dataIn2 = 32'd63; 
32'd1140: dataIn2 = 32'd56; 
32'd1141: dataIn2 = 32'd16; 
32'd1142: dataIn2 = 32'd44; 
32'd1143: dataIn2 = 32'd44; 
32'd1144: dataIn2 = 32'd87; 
32'd1145: dataIn2 = 32'd11; 
32'd1146: dataIn2 = 32'd0; 
32'd1147: dataIn2 = 32'd40; 
32'd1148: dataIn2 = 32'd22; 
32'd1149: dataIn2 = 32'd28; 
32'd1150: dataIn2 = 32'd77; 
32'd1151: dataIn2 = 32'd1; 
32'd1152: dataIn2 = 32'd24; 
32'd1153: dataIn2 = 32'd79; 
32'd1154: dataIn2 = 32'd5; 
32'd1155: dataIn2 = 32'd4; 
32'd1156: dataIn2 = 32'd77; 
32'd1157: dataIn2 = 32'd79; 
32'd1158: dataIn2 = 32'd38; 
32'd1159: dataIn2 = 32'd87; 
32'd1160: dataIn2 = 32'd73; 
32'd1161: dataIn2 = 32'd76; 
32'd1162: dataIn2 = 32'd64; 
32'd1163: dataIn2 = 32'd84; 
32'd1164: dataIn2 = 32'd29; 
32'd1165: dataIn2 = 32'd69; 
32'd1166: dataIn2 = 32'd74; 
32'd1167: dataIn2 = 32'd98; 
32'd1168: dataIn2 = 32'd92; 
32'd1169: dataIn2 = 32'd89; 
32'd1170: dataIn2 = 32'd44; 
32'd1171: dataIn2 = 32'd61; 
32'd1172: dataIn2 = 32'd78; 
32'd1173: dataIn2 = 32'd34; 
32'd1174: dataIn2 = 32'd66; 
32'd1175: dataIn2 = 32'd19; 
32'd1176: dataIn2 = 32'd21; 
32'd1177: dataIn2 = 32'd0; 
32'd1178: dataIn2 = 32'd15; 
32'd1179: dataIn2 = 32'd3; 
32'd1180: dataIn2 = 32'd72; 
32'd1181: dataIn2 = 32'd40; 
32'd1182: dataIn2 = 32'd26; 
32'd1183: dataIn2 = 32'd17; 
32'd1184: dataIn2 = 32'd60; 
32'd1185: dataIn2 = 32'd17; 
32'd1186: dataIn2 = 32'd8; 
32'd1187: dataIn2 = 32'd81; 
32'd1188: dataIn2 = 32'd85; 
32'd1189: dataIn2 = 32'd50; 
32'd1190: dataIn2 = 32'd100; 
32'd1191: dataIn2 = 32'd76; 
32'd1192: dataIn2 = 32'd48; 
32'd1193: dataIn2 = 32'd15; 
32'd1194: dataIn2 = 32'd70; 
32'd1195: dataIn2 = 32'd90; 
32'd1196: dataIn2 = 32'd2; 
32'd1197: dataIn2 = 32'd34; 
32'd1198: dataIn2 = 32'd31; 
32'd1199: dataIn2 = 32'd56; 
32'd1200: dataIn2 = 32'd68; 
32'd1201: dataIn2 = 32'd52; 
32'd1202: dataIn2 = 32'd79; 
32'd1203: dataIn2 = 32'd25; 
32'd1204: dataIn2 = 32'd17; 
32'd1205: dataIn2 = 32'd84; 
32'd1206: dataIn2 = 32'd83; 
32'd1207: dataIn2 = 32'd89; 
32'd1208: dataIn2 = 32'd63; 
32'd1209: dataIn2 = 32'd77; 
32'd1210: dataIn2 = 32'd56; 
32'd1211: dataIn2 = 32'd0; 
32'd1212: dataIn2 = 32'd18; 
32'd1213: dataIn2 = 32'd84; 
32'd1214: dataIn2 = 32'd5; 
32'd1215: dataIn2 = 32'd23; 
32'd1216: dataIn2 = 32'd34; 
32'd1217: dataIn2 = 32'd71; 
32'd1218: dataIn2 = 32'd64; 
32'd1219: dataIn2 = 32'd72; 
32'd1220: dataIn2 = 32'd63; 
32'd1221: dataIn2 = 32'd15; 
32'd1222: dataIn2 = 32'd67; 
32'd1223: dataIn2 = 32'd41; 
32'd1224: dataIn2 = 32'd100; 
32'd1225: dataIn2 = 32'd16; 
32'd1226: dataIn2 = 32'd2; 
32'd1227: dataIn2 = 32'd76; 
32'd1228: dataIn2 = 32'd54; 
32'd1229: dataIn2 = 32'd0; 
32'd1230: dataIn2 = 32'd76; 
32'd1231: dataIn2 = 32'd53; 
32'd1232: dataIn2 = 32'd24; 
32'd1233: dataIn2 = 32'd83; 
32'd1234: dataIn2 = 32'd22; 
32'd1235: dataIn2 = 32'd68; 
32'd1236: dataIn2 = 32'd95; 
32'd1237: dataIn2 = 32'd18; 
32'd1238: dataIn2 = 32'd100; 
32'd1239: dataIn2 = 32'd75; 
32'd1240: dataIn2 = 32'd30; 
32'd1241: dataIn2 = 32'd88; 
32'd1242: dataIn2 = 32'd7; 
32'd1243: dataIn2 = 32'd94; 
32'd1244: dataIn2 = 32'd61; 
32'd1245: dataIn2 = 32'd73; 
32'd1246: dataIn2 = 32'd42; 
32'd1247: dataIn2 = 32'd33; 
32'd1248: dataIn2 = 32'd13; 
32'd1249: dataIn2 = 32'd9; 
32'd1250: dataIn2 = 32'd91; 
32'd1251: dataIn2 = 32'd100; 
32'd1252: dataIn2 = 32'd12; 
32'd1253: dataIn2 = 32'd13; 
32'd1254: dataIn2 = 32'd64; 
32'd1255: dataIn2 = 32'd33; 
32'd1256: dataIn2 = 32'd90; 
32'd1257: dataIn2 = 32'd100; 
32'd1258: dataIn2 = 32'd60; 
32'd1259: dataIn2 = 32'd51; 
32'd1260: dataIn2 = 32'd68; 
32'd1261: dataIn2 = 32'd44; 
32'd1262: dataIn2 = 32'd56; 
32'd1263: dataIn2 = 32'd66; 
32'd1264: dataIn2 = 32'd5; 
32'd1265: dataIn2 = 32'd43; 
32'd1266: dataIn2 = 32'd42; 
32'd1267: dataIn2 = 32'd40; 
32'd1268: dataIn2 = 32'd42; 
32'd1269: dataIn2 = 32'd56; 
32'd1270: dataIn2 = 32'd71; 
32'd1271: dataIn2 = 32'd13; 
32'd1272: dataIn2 = 32'd14; 
32'd1273: dataIn2 = 32'd74; 
32'd1274: dataIn2 = 32'd96; 
32'd1275: dataIn2 = 32'd80; 
32'd1276: dataIn2 = 32'd79; 
32'd1277: dataIn2 = 32'd35; 
32'd1278: dataIn2 = 32'd40; 
32'd1279: dataIn2 = 32'd3; 
32'd1280: dataIn2 = 32'd16; 
32'd1281: dataIn2 = 32'd99; 
32'd1282: dataIn2 = 32'd34; 
32'd1283: dataIn2 = 32'd38; 
32'd1284: dataIn2 = 32'd69; 
32'd1285: dataIn2 = 32'd90; 
32'd1286: dataIn2 = 32'd74; 
32'd1287: dataIn2 = 32'd64; 
32'd1288: dataIn2 = 32'd49; 
32'd1289: dataIn2 = 32'd70; 
32'd1290: dataIn2 = 32'd19; 
32'd1291: dataIn2 = 32'd46; 
32'd1292: dataIn2 = 32'd7; 
32'd1293: dataIn2 = 32'd54; 
32'd1294: dataIn2 = 32'd91; 
32'd1295: dataIn2 = 32'd24; 
32'd1296: dataIn2 = 32'd12; 
32'd1297: dataIn2 = 32'd9; 
32'd1298: dataIn2 = 32'd95; 
32'd1299: dataIn2 = 32'd87; 
32'd1300: dataIn2 = 32'd52; 
32'd1301: dataIn2 = 32'd16; 
32'd1302: dataIn2 = 32'd81; 
32'd1303: dataIn2 = 32'd91; 
32'd1304: dataIn2 = 32'd38; 
32'd1305: dataIn2 = 32'd44; 
32'd1306: dataIn2 = 32'd4; 
32'd1307: dataIn2 = 32'd62; 
32'd1308: dataIn2 = 32'd18; 
32'd1309: dataIn2 = 32'd63; 
32'd1310: dataIn2 = 32'd50; 
32'd1311: dataIn2 = 32'd14; 
32'd1312: dataIn2 = 32'd79; 
32'd1313: dataIn2 = 32'd67; 
32'd1314: dataIn2 = 32'd78; 
32'd1315: dataIn2 = 32'd53; 
32'd1316: dataIn2 = 32'd3; 
32'd1317: dataIn2 = 32'd47; 
32'd1318: dataIn2 = 32'd15; 
32'd1319: dataIn2 = 32'd20; 
32'd1320: dataIn2 = 32'd18; 
32'd1321: dataIn2 = 32'd51; 
32'd1322: dataIn2 = 32'd17; 
32'd1323: dataIn2 = 32'd68; 
32'd1324: dataIn2 = 32'd54; 
32'd1325: dataIn2 = 32'd82; 
32'd1326: dataIn2 = 32'd48; 
32'd1327: dataIn2 = 32'd93; 
32'd1328: dataIn2 = 32'd68; 
32'd1329: dataIn2 = 32'd20; 
32'd1330: dataIn2 = 32'd98; 
32'd1331: dataIn2 = 32'd67; 
32'd1332: dataIn2 = 32'd97; 
32'd1333: dataIn2 = 32'd19; 
32'd1334: dataIn2 = 32'd3; 
32'd1335: dataIn2 = 32'd35; 
32'd1336: dataIn2 = 32'd42; 
32'd1337: dataIn2 = 32'd92; 
32'd1338: dataIn2 = 32'd67; 
32'd1339: dataIn2 = 32'd13; 
32'd1340: dataIn2 = 32'd74; 
32'd1341: dataIn2 = 32'd100; 
32'd1342: dataIn2 = 32'd29; 
32'd1343: dataIn2 = 32'd45; 
32'd1344: dataIn2 = 32'd60; 
32'd1345: dataIn2 = 32'd24; 
32'd1346: dataIn2 = 32'd55; 
32'd1347: dataIn2 = 32'd61; 
32'd1348: dataIn2 = 32'd29; 
32'd1349: dataIn2 = 32'd9; 
32'd1350: dataIn2 = 32'd45; 
32'd1351: dataIn2 = 32'd16; 
32'd1352: dataIn2 = 32'd90; 
32'd1353: dataIn2 = 32'd59; 
32'd1354: dataIn2 = 32'd34; 
32'd1355: dataIn2 = 32'd32; 
32'd1356: dataIn2 = 32'd63; 
32'd1357: dataIn2 = 32'd5; 
32'd1358: dataIn2 = 32'd4; 
32'd1359: dataIn2 = 32'd93; 
32'd1360: dataIn2 = 32'd88; 
32'd1361: dataIn2 = 32'd83; 
32'd1362: dataIn2 = 32'd57; 
32'd1363: dataIn2 = 32'd68; 
32'd1364: dataIn2 = 32'd68; 
32'd1365: dataIn2 = 32'd85; 
32'd1366: dataIn2 = 32'd22; 
32'd1367: dataIn2 = 32'd0; 
32'd1368: dataIn2 = 32'd18; 
32'd1369: dataIn2 = 32'd26; 
32'd1370: dataIn2 = 32'd33; 
32'd1371: dataIn2 = 32'd38; 
32'd1372: dataIn2 = 32'd92; 
32'd1373: dataIn2 = 32'd48; 
32'd1374: dataIn2 = 32'd94; 
32'd1375: dataIn2 = 32'd45; 
32'd1376: dataIn2 = 32'd30; 
32'd1377: dataIn2 = 32'd42; 
32'd1378: dataIn2 = 32'd9; 
32'd1379: dataIn2 = 32'd10; 
32'd1380: dataIn2 = 32'd57; 
32'd1381: dataIn2 = 32'd7; 
32'd1382: dataIn2 = 32'd13; 
32'd1383: dataIn2 = 32'd30; 
32'd1384: dataIn2 = 32'd37; 
32'd1385: dataIn2 = 32'd65; 
32'd1386: dataIn2 = 32'd54; 
32'd1387: dataIn2 = 32'd22; 
32'd1388: dataIn2 = 32'd92; 
32'd1389: dataIn2 = 32'd72; 
32'd1390: dataIn2 = 32'd34; 
32'd1391: dataIn2 = 32'd43; 
32'd1392: dataIn2 = 32'd29; 
32'd1393: dataIn2 = 32'd53; 
32'd1394: dataIn2 = 32'd22; 
32'd1395: dataIn2 = 32'd48; 
32'd1396: dataIn2 = 32'd58; 
32'd1397: dataIn2 = 32'd57; 
32'd1398: dataIn2 = 32'd44; 
32'd1399: dataIn2 = 32'd74; 
32'd1400: dataIn2 = 32'd6; 
32'd1401: dataIn2 = 32'd6; 
32'd1402: dataIn2 = 32'd49; 
32'd1403: dataIn2 = 32'd62; 
32'd1404: dataIn2 = 32'd11; 
32'd1405: dataIn2 = 32'd64; 
32'd1406: dataIn2 = 32'd97; 
32'd1407: dataIn2 = 32'd74; 
32'd1408: dataIn2 = 32'd50; 
32'd1409: dataIn2 = 32'd19; 
32'd1410: dataIn2 = 32'd92; 
32'd1411: dataIn2 = 32'd21; 
32'd1412: dataIn2 = 32'd53; 
32'd1413: dataIn2 = 32'd64; 
32'd1414: dataIn2 = 32'd46; 
32'd1415: dataIn2 = 32'd39; 
32'd1416: dataIn2 = 32'd10; 
32'd1417: dataIn2 = 32'd25; 
32'd1418: dataIn2 = 32'd32; 
32'd1419: dataIn2 = 32'd37; 
32'd1420: dataIn2 = 32'd9; 
32'd1421: dataIn2 = 32'd61; 
32'd1422: dataIn2 = 32'd25; 
32'd1423: dataIn2 = 32'd38; 
32'd1424: dataIn2 = 32'd27; 
32'd1425: dataIn2 = 32'd13; 
32'd1426: dataIn2 = 32'd44; 
32'd1427: dataIn2 = 32'd51; 
32'd1428: dataIn2 = 32'd5; 
32'd1429: dataIn2 = 32'd86; 
32'd1430: dataIn2 = 32'd91; 
32'd1431: dataIn2 = 32'd14; 
32'd1432: dataIn2 = 32'd87; 
32'd1433: dataIn2 = 32'd96; 
32'd1434: dataIn2 = 32'd59; 
32'd1435: dataIn2 = 32'd51; 
32'd1436: dataIn2 = 32'd28; 
32'd1437: dataIn2 = 32'd4; 
32'd1438: dataIn2 = 32'd27; 
32'd1439: dataIn2 = 32'd77; 
32'd1440: dataIn2 = 32'd21; 
32'd1441: dataIn2 = 32'd34; 
32'd1442: dataIn2 = 32'd88; 
32'd1443: dataIn2 = 32'd12; 
32'd1444: dataIn2 = 32'd0; 
32'd1445: dataIn2 = 32'd19; 
32'd1446: dataIn2 = 32'd29; 
32'd1447: dataIn2 = 32'd2; 
32'd1448: dataIn2 = 32'd19; 
32'd1449: dataIn2 = 32'd57; 
32'd1450: dataIn2 = 32'd86; 
32'd1451: dataIn2 = 32'd89; 
32'd1452: dataIn2 = 32'd97; 
32'd1453: dataIn2 = 32'd5; 
32'd1454: dataIn2 = 32'd8; 
32'd1455: dataIn2 = 32'd49; 
32'd1456: dataIn2 = 32'd49; 
32'd1457: dataIn2 = 32'd93; 
32'd1458: dataIn2 = 32'd66; 
32'd1459: dataIn2 = 32'd50; 
32'd1460: dataIn2 = 32'd65; 
32'd1461: dataIn2 = 32'd93; 
32'd1462: dataIn2 = 32'd62; 
32'd1463: dataIn2 = 32'd93; 
32'd1464: dataIn2 = 32'd83; 
32'd1465: dataIn2 = 32'd93; 
32'd1466: dataIn2 = 32'd69; 
32'd1467: dataIn2 = 32'd44; 
32'd1468: dataIn2 = 32'd76; 
32'd1469: dataIn2 = 32'd2; 
32'd1470: dataIn2 = 32'd4; 
32'd1471: dataIn2 = 32'd52; 
32'd1472: dataIn2 = 32'd96; 
32'd1473: dataIn2 = 32'd47; 
32'd1474: dataIn2 = 32'd96; 
32'd1475: dataIn2 = 32'd73; 
32'd1476: dataIn2 = 32'd96; 
32'd1477: dataIn2 = 32'd80; 
32'd1478: dataIn2 = 32'd59; 
32'd1479: dataIn2 = 32'd2; 
32'd1480: dataIn2 = 32'd37; 
32'd1481: dataIn2 = 32'd92; 
32'd1482: dataIn2 = 32'd54; 
32'd1483: dataIn2 = 32'd83; 
32'd1484: dataIn2 = 32'd48; 
32'd1485: dataIn2 = 32'd1; 
32'd1486: dataIn2 = 32'd76; 
32'd1487: dataIn2 = 32'd90; 
32'd1488: dataIn2 = 32'd17; 
32'd1489: dataIn2 = 32'd76; 
32'd1490: dataIn2 = 32'd79; 
32'd1491: dataIn2 = 32'd92; 
32'd1492: dataIn2 = 32'd61; 
32'd1493: dataIn2 = 32'd30; 
32'd1494: dataIn2 = 32'd1; 
32'd1495: dataIn2 = 32'd6; 
32'd1496: dataIn2 = 32'd84; 
32'd1497: dataIn2 = 32'd40; 
32'd1498: dataIn2 = 32'd47; 
32'd1499: dataIn2 = 32'd11; 
32'd1500: dataIn2 = 32'd91; 
32'd1501: dataIn2 = 32'd46; 
32'd1502: dataIn2 = 32'd4; 
32'd1503: dataIn2 = 32'd58; 
32'd1504: dataIn2 = 32'd38; 
32'd1505: dataIn2 = 32'd70; 
32'd1506: dataIn2 = 32'd17; 
32'd1507: dataIn2 = 32'd6; 
32'd1508: dataIn2 = 32'd14; 
32'd1509: dataIn2 = 32'd42; 
32'd1510: dataIn2 = 32'd84; 
32'd1511: dataIn2 = 32'd48; 
32'd1512: dataIn2 = 32'd35; 
32'd1513: dataIn2 = 32'd28; 
32'd1514: dataIn2 = 32'd14; 
32'd1515: dataIn2 = 32'd75; 
32'd1516: dataIn2 = 32'd40; 
32'd1517: dataIn2 = 32'd20; 
32'd1518: dataIn2 = 32'd56; 
32'd1519: dataIn2 = 32'd24; 
32'd1520: dataIn2 = 32'd42; 
32'd1521: dataIn2 = 32'd81; 
32'd1522: dataIn2 = 32'd24; 
32'd1523: dataIn2 = 32'd26; 
32'd1524: dataIn2 = 32'd13; 
32'd1525: dataIn2 = 32'd89; 
32'd1526: dataIn2 = 32'd37; 
32'd1527: dataIn2 = 32'd68; 
32'd1528: dataIn2 = 32'd69; 
32'd1529: dataIn2 = 32'd19; 
32'd1530: dataIn2 = 32'd67; 
32'd1531: dataIn2 = 32'd9; 
32'd1532: dataIn2 = 32'd38; 
32'd1533: dataIn2 = 32'd19; 
32'd1534: dataIn2 = 32'd67; 
32'd1535: dataIn2 = 32'd58; 
32'd1536: dataIn2 = 32'd31; 
32'd1537: dataIn2 = 32'd56; 
32'd1538: dataIn2 = 32'd38; 
32'd1539: dataIn2 = 32'd89; 
32'd1540: dataIn2 = 32'd80; 
32'd1541: dataIn2 = 32'd54; 
32'd1542: dataIn2 = 32'd51; 
32'd1543: dataIn2 = 32'd47; 
32'd1544: dataIn2 = 32'd61; 
32'd1545: dataIn2 = 32'd82; 
32'd1546: dataIn2 = 32'd0; 
32'd1547: dataIn2 = 32'd100; 
32'd1548: dataIn2 = 32'd11; 
32'd1549: dataIn2 = 32'd85; 
32'd1550: dataIn2 = 32'd64; 
32'd1551: dataIn2 = 32'd65; 
32'd1552: dataIn2 = 32'd7; 
32'd1553: dataIn2 = 32'd41; 
32'd1554: dataIn2 = 32'd95; 
32'd1555: dataIn2 = 32'd0; 
32'd1556: dataIn2 = 32'd8; 
32'd1557: dataIn2 = 32'd15; 
32'd1558: dataIn2 = 32'd60; 
32'd1559: dataIn2 = 32'd49; 
32'd1560: dataIn2 = 32'd0; 
32'd1561: dataIn2 = 32'd84; 
32'd1562: dataIn2 = 32'd52; 
32'd1563: dataIn2 = 32'd42; 
32'd1564: dataIn2 = 32'd36; 
32'd1565: dataIn2 = 32'd49; 
32'd1566: dataIn2 = 32'd22; 
32'd1567: dataIn2 = 32'd46; 
32'd1568: dataIn2 = 32'd4; 
32'd1569: dataIn2 = 32'd74; 
32'd1570: dataIn2 = 32'd6; 
32'd1571: dataIn2 = 32'd42; 
32'd1572: dataIn2 = 32'd3; 
32'd1573: dataIn2 = 32'd13; 
32'd1574: dataIn2 = 32'd25; 
32'd1575: dataIn2 = 32'd1; 
32'd1576: dataIn2 = 32'd17; 
32'd1577: dataIn2 = 32'd94; 
32'd1578: dataIn2 = 32'd6; 
32'd1579: dataIn2 = 32'd46; 
32'd1580: dataIn2 = 32'd25; 
32'd1581: dataIn2 = 32'd11; 
32'd1582: dataIn2 = 32'd62; 
32'd1583: dataIn2 = 32'd77; 
32'd1584: dataIn2 = 32'd88; 
32'd1585: dataIn2 = 32'd53; 
32'd1586: dataIn2 = 32'd69; 
32'd1587: dataIn2 = 32'd8; 
32'd1588: dataIn2 = 32'd93; 
32'd1589: dataIn2 = 32'd26; 
32'd1590: dataIn2 = 32'd44; 
32'd1591: dataIn2 = 32'd12; 
32'd1592: dataIn2 = 32'd83; 
32'd1593: dataIn2 = 32'd5; 
32'd1594: dataIn2 = 32'd96; 
32'd1595: dataIn2 = 32'd6; 
32'd1596: dataIn2 = 32'd63; 
32'd1597: dataIn2 = 32'd88; 
32'd1598: dataIn2 = 32'd0; 
32'd1599: dataIn2 = 32'd79; 
32'd1600: dataIn2 = 32'd91; 
32'd1601: dataIn2 = 32'd85; 
32'd1602: dataIn2 = 32'd37; 
32'd1603: dataIn2 = 32'd1; 
32'd1604: dataIn2 = 32'd79; 
32'd1605: dataIn2 = 32'd40; 
32'd1606: dataIn2 = 32'd51; 
32'd1607: dataIn2 = 32'd50; 
32'd1608: dataIn2 = 32'd50; 
32'd1609: dataIn2 = 32'd34; 
32'd1610: dataIn2 = 32'd53; 
32'd1611: dataIn2 = 32'd46; 
32'd1612: dataIn2 = 32'd33; 
32'd1613: dataIn2 = 32'd25; 
32'd1614: dataIn2 = 32'd48; 
32'd1615: dataIn2 = 32'd84; 
32'd1616: dataIn2 = 32'd59; 
32'd1617: dataIn2 = 32'd26; 
32'd1618: dataIn2 = 32'd82; 
32'd1619: dataIn2 = 32'd37; 
32'd1620: dataIn2 = 32'd89; 
32'd1621: dataIn2 = 32'd51; 
32'd1622: dataIn2 = 32'd95; 
32'd1623: dataIn2 = 32'd58; 
32'd1624: dataIn2 = 32'd11; 
32'd1625: dataIn2 = 32'd8; 
32'd1626: dataIn2 = 32'd98; 
32'd1627: dataIn2 = 32'd21; 
32'd1628: dataIn2 = 32'd57; 
32'd1629: dataIn2 = 32'd65; 
32'd1630: dataIn2 = 32'd1; 
32'd1631: dataIn2 = 32'd79; 
32'd1632: dataIn2 = 32'd93; 
32'd1633: dataIn2 = 32'd17; 
32'd1634: dataIn2 = 32'd21; 
32'd1635: dataIn2 = 32'd6; 
32'd1636: dataIn2 = 32'd11; 
32'd1637: dataIn2 = 32'd46; 
32'd1638: dataIn2 = 32'd93; 
32'd1639: dataIn2 = 32'd80; 
32'd1640: dataIn2 = 32'd43; 
32'd1641: dataIn2 = 32'd33; 
32'd1642: dataIn2 = 32'd20; 
32'd1643: dataIn2 = 32'd8; 
32'd1644: dataIn2 = 32'd51; 
32'd1645: dataIn2 = 32'd74; 
32'd1646: dataIn2 = 32'd37; 
32'd1647: dataIn2 = 32'd64; 
32'd1648: dataIn2 = 32'd36; 
32'd1649: dataIn2 = 32'd73; 
32'd1650: dataIn2 = 32'd51; 
32'd1651: dataIn2 = 32'd75; 
32'd1652: dataIn2 = 32'd48; 
32'd1653: dataIn2 = 32'd72; 
32'd1654: dataIn2 = 32'd2; 
32'd1655: dataIn2 = 32'd64; 
32'd1656: dataIn2 = 32'd54; 
32'd1657: dataIn2 = 32'd66; 
32'd1658: dataIn2 = 32'd31; 
32'd1659: dataIn2 = 32'd84; 
32'd1660: dataIn2 = 32'd76; 
32'd1661: dataIn2 = 32'd24; 
32'd1662: dataIn2 = 32'd40; 
32'd1663: dataIn2 = 32'd33; 
32'd1664: dataIn2 = 32'd57; 
32'd1665: dataIn2 = 32'd55; 
32'd1666: dataIn2 = 32'd55; 
32'd1667: dataIn2 = 32'd19; 
32'd1668: dataIn2 = 32'd84; 
32'd1669: dataIn2 = 32'd27; 
32'd1670: dataIn2 = 32'd52; 
32'd1671: dataIn2 = 32'd62; 
32'd1672: dataIn2 = 32'd41; 
32'd1673: dataIn2 = 32'd14; 
32'd1674: dataIn2 = 32'd97; 
32'd1675: dataIn2 = 32'd32; 
32'd1676: dataIn2 = 32'd49; 
32'd1677: dataIn2 = 32'd94; 
32'd1678: dataIn2 = 32'd23; 
32'd1679: dataIn2 = 32'd28; 
32'd1680: dataIn2 = 32'd5; 
32'd1681: dataIn2 = 32'd15; 
32'd1682: dataIn2 = 32'd19; 
32'd1683: dataIn2 = 32'd68; 
32'd1684: dataIn2 = 32'd2; 
32'd1685: dataIn2 = 32'd98; 
32'd1686: dataIn2 = 32'd19; 
32'd1687: dataIn2 = 32'd59; 
32'd1688: dataIn2 = 32'd40; 
32'd1689: dataIn2 = 32'd75; 
32'd1690: dataIn2 = 32'd26; 
32'd1691: dataIn2 = 32'd13; 
32'd1692: dataIn2 = 32'd52; 
32'd1693: dataIn2 = 32'd86; 
32'd1694: dataIn2 = 32'd6; 
32'd1695: dataIn2 = 32'd65; 
32'd1696: dataIn2 = 32'd80; 
32'd1697: dataIn2 = 32'd26; 
32'd1698: dataIn2 = 32'd62; 
32'd1699: dataIn2 = 32'd81; 
32'd1700: dataIn2 = 32'd57; 
32'd1701: dataIn2 = 32'd0; 
32'd1702: dataIn2 = 32'd50; 
32'd1703: dataIn2 = 32'd53; 
32'd1704: dataIn2 = 32'd7; 
32'd1705: dataIn2 = 32'd94; 
32'd1706: dataIn2 = 32'd52; 
32'd1707: dataIn2 = 32'd7; 
32'd1708: dataIn2 = 32'd60; 
32'd1709: dataIn2 = 32'd3; 
32'd1710: dataIn2 = 32'd87; 
32'd1711: dataIn2 = 32'd71; 
32'd1712: dataIn2 = 32'd8; 
32'd1713: dataIn2 = 32'd3; 
32'd1714: dataIn2 = 32'd75; 
32'd1715: dataIn2 = 32'd22; 
32'd1716: dataIn2 = 32'd17; 
32'd1717: dataIn2 = 32'd65; 
32'd1718: dataIn2 = 32'd65; 
32'd1719: dataIn2 = 32'd81; 
32'd1720: dataIn2 = 32'd72; 
32'd1721: dataIn2 = 32'd76; 
32'd1722: dataIn2 = 32'd64; 
32'd1723: dataIn2 = 32'd88; 
32'd1724: dataIn2 = 32'd19; 
32'd1725: dataIn2 = 32'd95; 
32'd1726: dataIn2 = 32'd38; 
32'd1727: dataIn2 = 32'd75; 
32'd1728: dataIn2 = 32'd59; 
32'd1729: dataIn2 = 32'd31; 
32'd1730: dataIn2 = 32'd17; 
32'd1731: dataIn2 = 32'd7; 
32'd1732: dataIn2 = 32'd55; 
32'd1733: dataIn2 = 32'd44; 
32'd1734: dataIn2 = 32'd39; 
32'd1735: dataIn2 = 32'd73; 
32'd1736: dataIn2 = 32'd0; 
32'd1737: dataIn2 = 32'd57; 
32'd1738: dataIn2 = 32'd27; 
32'd1739: dataIn2 = 32'd71; 
32'd1740: dataIn2 = 32'd87; 
32'd1741: dataIn2 = 32'd65; 
32'd1742: dataIn2 = 32'd31; 
32'd1743: dataIn2 = 32'd100; 
32'd1744: dataIn2 = 32'd40; 
32'd1745: dataIn2 = 32'd86; 
32'd1746: dataIn2 = 32'd8; 
32'd1747: dataIn2 = 32'd75; 
32'd1748: dataIn2 = 32'd35; 
32'd1749: dataIn2 = 32'd53; 
32'd1750: dataIn2 = 32'd100; 
32'd1751: dataIn2 = 32'd14; 
32'd1752: dataIn2 = 32'd95; 
32'd1753: dataIn2 = 32'd88; 
32'd1754: dataIn2 = 32'd89; 
32'd1755: dataIn2 = 32'd9; 
32'd1756: dataIn2 = 32'd80; 
32'd1757: dataIn2 = 32'd55; 
32'd1758: dataIn2 = 32'd14; 
32'd1759: dataIn2 = 32'd33; 
32'd1760: dataIn2 = 32'd93; 
32'd1761: dataIn2 = 32'd91; 
32'd1762: dataIn2 = 32'd58; 
32'd1763: dataIn2 = 32'd88; 
32'd1764: dataIn2 = 32'd6; 
32'd1765: dataIn2 = 32'd46; 
32'd1766: dataIn2 = 32'd14; 
32'd1767: dataIn2 = 32'd25; 
32'd1768: dataIn2 = 32'd69; 
32'd1769: dataIn2 = 32'd61; 
32'd1770: dataIn2 = 32'd81; 
32'd1771: dataIn2 = 32'd6; 
32'd1772: dataIn2 = 32'd88; 
32'd1773: dataIn2 = 32'd48; 
32'd1774: dataIn2 = 32'd45; 
32'd1775: dataIn2 = 32'd83; 
32'd1776: dataIn2 = 32'd58; 
32'd1777: dataIn2 = 32'd85; 
32'd1778: dataIn2 = 32'd57; 
32'd1779: dataIn2 = 32'd17; 
32'd1780: dataIn2 = 32'd5; 
32'd1781: dataIn2 = 32'd58; 
32'd1782: dataIn2 = 32'd29; 
32'd1783: dataIn2 = 32'd17; 
32'd1784: dataIn2 = 32'd86; 
32'd1785: dataIn2 = 32'd13; 
32'd1786: dataIn2 = 32'd29; 
32'd1787: dataIn2 = 32'd34; 
32'd1788: dataIn2 = 32'd14; 
32'd1789: dataIn2 = 32'd38; 
32'd1790: dataIn2 = 32'd46; 
32'd1791: dataIn2 = 32'd17; 
32'd1792: dataIn2 = 32'd74; 
32'd1793: dataIn2 = 32'd79; 
32'd1794: dataIn2 = 32'd46; 
32'd1795: dataIn2 = 32'd28; 
32'd1796: dataIn2 = 32'd73; 
32'd1797: dataIn2 = 32'd84; 
32'd1798: dataIn2 = 32'd82; 
32'd1799: dataIn2 = 32'd65; 
32'd1800: dataIn2 = 32'd7; 
32'd1801: dataIn2 = 32'd13; 
32'd1802: dataIn2 = 32'd83; 
32'd1803: dataIn2 = 32'd86; 
32'd1804: dataIn2 = 32'd38; 
32'd1805: dataIn2 = 32'd88; 
32'd1806: dataIn2 = 32'd94; 
32'd1807: dataIn2 = 32'd52; 
32'd1808: dataIn2 = 32'd63; 
32'd1809: dataIn2 = 32'd22; 
32'd1810: dataIn2 = 32'd84; 
32'd1811: dataIn2 = 32'd95; 
32'd1812: dataIn2 = 32'd65; 
32'd1813: dataIn2 = 32'd49; 
32'd1814: dataIn2 = 32'd0; 
32'd1815: dataIn2 = 32'd87; 
32'd1816: dataIn2 = 32'd53; 
32'd1817: dataIn2 = 32'd29; 
32'd1818: dataIn2 = 32'd28; 
32'd1819: dataIn2 = 32'd19; 
32'd1820: dataIn2 = 32'd53; 
32'd1821: dataIn2 = 32'd86; 
32'd1822: dataIn2 = 32'd12; 
32'd1823: dataIn2 = 32'd46; 
32'd1824: dataIn2 = 32'd2; 
32'd1825: dataIn2 = 32'd35; 
32'd1826: dataIn2 = 32'd31; 
32'd1827: dataIn2 = 32'd28; 
32'd1828: dataIn2 = 32'd4; 
32'd1829: dataIn2 = 32'd94; 
32'd1830: dataIn2 = 32'd45; 
32'd1831: dataIn2 = 32'd80; 
32'd1832: dataIn2 = 32'd75; 
32'd1833: dataIn2 = 32'd20; 
32'd1834: dataIn2 = 32'd61; 
32'd1835: dataIn2 = 32'd15; 
32'd1836: dataIn2 = 32'd62; 
32'd1837: dataIn2 = 32'd18; 
32'd1838: dataIn2 = 32'd50; 
32'd1839: dataIn2 = 32'd19; 
32'd1840: dataIn2 = 32'd78; 
32'd1841: dataIn2 = 32'd74; 
32'd1842: dataIn2 = 32'd39; 
32'd1843: dataIn2 = 32'd12; 
32'd1844: dataIn2 = 32'd22; 
32'd1845: dataIn2 = 32'd68; 
32'd1846: dataIn2 = 32'd69; 
32'd1847: dataIn2 = 32'd27; 
32'd1848: dataIn2 = 32'd72; 
32'd1849: dataIn2 = 32'd63; 
32'd1850: dataIn2 = 32'd39; 
32'd1851: dataIn2 = 32'd4; 
32'd1852: dataIn2 = 32'd20; 
32'd1853: dataIn2 = 32'd2; 
32'd1854: dataIn2 = 32'd0; 
32'd1855: dataIn2 = 32'd80; 
32'd1856: dataIn2 = 32'd91; 
32'd1857: dataIn2 = 32'd47; 
32'd1858: dataIn2 = 32'd27; 
32'd1859: dataIn2 = 32'd16; 
32'd1860: dataIn2 = 32'd77; 
32'd1861: dataIn2 = 32'd48; 
32'd1862: dataIn2 = 32'd52; 
32'd1863: dataIn2 = 32'd14; 
32'd1864: dataIn2 = 32'd14; 
32'd1865: dataIn2 = 32'd67; 
32'd1866: dataIn2 = 32'd51; 
32'd1867: dataIn2 = 32'd96; 
32'd1868: dataIn2 = 32'd59; 
32'd1869: dataIn2 = 32'd33; 
32'd1870: dataIn2 = 32'd45; 
32'd1871: dataIn2 = 32'd11; 
32'd1872: dataIn2 = 32'd64; 
32'd1873: dataIn2 = 32'd99; 
32'd1874: dataIn2 = 32'd30; 
32'd1875: dataIn2 = 32'd41; 
32'd1876: dataIn2 = 32'd36; 
32'd1877: dataIn2 = 32'd28; 
32'd1878: dataIn2 = 32'd58; 
32'd1879: dataIn2 = 32'd1; 
32'd1880: dataIn2 = 32'd7; 
32'd1881: dataIn2 = 32'd80; 
32'd1882: dataIn2 = 32'd31; 
32'd1883: dataIn2 = 32'd80; 
32'd1884: dataIn2 = 32'd75; 
32'd1885: dataIn2 = 32'd76; 
32'd1886: dataIn2 = 32'd91; 
32'd1887: dataIn2 = 32'd1; 
32'd1888: dataIn2 = 32'd0; 
32'd1889: dataIn2 = 32'd53; 
32'd1890: dataIn2 = 32'd45; 
32'd1891: dataIn2 = 32'd96; 
32'd1892: dataIn2 = 32'd51; 
32'd1893: dataIn2 = 32'd62; 
32'd1894: dataIn2 = 32'd31; 
32'd1895: dataIn2 = 32'd85; 
32'd1896: dataIn2 = 32'd98; 
32'd1897: dataIn2 = 32'd100; 
32'd1898: dataIn2 = 32'd91; 
32'd1899: dataIn2 = 32'd93; 
32'd1900: dataIn2 = 32'd27; 
32'd1901: dataIn2 = 32'd10; 
32'd1902: dataIn2 = 32'd34; 
32'd1903: dataIn2 = 32'd61; 
32'd1904: dataIn2 = 32'd24; 
32'd1905: dataIn2 = 32'd8; 
32'd1906: dataIn2 = 32'd80; 
32'd1907: dataIn2 = 32'd93; 
32'd1908: dataIn2 = 32'd34; 
32'd1909: dataIn2 = 32'd22; 
32'd1910: dataIn2 = 32'd45; 
32'd1911: dataIn2 = 32'd46; 
32'd1912: dataIn2 = 32'd30; 
32'd1913: dataIn2 = 32'd37; 
32'd1914: dataIn2 = 32'd95; 
32'd1915: dataIn2 = 32'd17; 
32'd1916: dataIn2 = 32'd33; 
32'd1917: dataIn2 = 32'd58; 
32'd1918: dataIn2 = 32'd84; 
32'd1919: dataIn2 = 32'd16; 
32'd1920: dataIn2 = 32'd82; 
32'd1921: dataIn2 = 32'd79; 
32'd1922: dataIn2 = 32'd71; 
32'd1923: dataIn2 = 32'd55; 
32'd1924: dataIn2 = 32'd2; 
32'd1925: dataIn2 = 32'd4; 
32'd1926: dataIn2 = 32'd96; 
32'd1927: dataIn2 = 32'd22; 
32'd1928: dataIn2 = 32'd10; 
32'd1929: dataIn2 = 32'd58; 
32'd1930: dataIn2 = 32'd19; 
32'd1931: dataIn2 = 32'd46; 
32'd1932: dataIn2 = 32'd27; 
32'd1933: dataIn2 = 32'd39; 
32'd1934: dataIn2 = 32'd30; 
32'd1935: dataIn2 = 32'd38; 
32'd1936: dataIn2 = 32'd56; 
32'd1937: dataIn2 = 32'd85; 
32'd1938: dataIn2 = 32'd30; 
32'd1939: dataIn2 = 32'd64; 
32'd1940: dataIn2 = 32'd44; 
32'd1941: dataIn2 = 32'd13; 
32'd1942: dataIn2 = 32'd96; 
32'd1943: dataIn2 = 32'd37; 
32'd1944: dataIn2 = 32'd35; 
32'd1945: dataIn2 = 32'd93; 
32'd1946: dataIn2 = 32'd2; 
32'd1947: dataIn2 = 32'd39; 
32'd1948: dataIn2 = 32'd44; 
32'd1949: dataIn2 = 32'd11; 
32'd1950: dataIn2 = 32'd60; 
32'd1951: dataIn2 = 32'd8; 
32'd1952: dataIn2 = 32'd41; 
32'd1953: dataIn2 = 32'd90; 
32'd1954: dataIn2 = 32'd26; 
32'd1955: dataIn2 = 32'd8; 
32'd1956: dataIn2 = 32'd85; 
32'd1957: dataIn2 = 32'd25; 
32'd1958: dataIn2 = 32'd45; 
32'd1959: dataIn2 = 32'd65; 
32'd1960: dataIn2 = 32'd34; 
32'd1961: dataIn2 = 32'd84; 
32'd1962: dataIn2 = 32'd22; 
32'd1963: dataIn2 = 32'd80; 
32'd1964: dataIn2 = 32'd47; 
32'd1965: dataIn2 = 32'd79; 
32'd1966: dataIn2 = 32'd54; 
32'd1967: dataIn2 = 32'd36; 
32'd1968: dataIn2 = 32'd89; 
32'd1969: dataIn2 = 32'd35; 
32'd1970: dataIn2 = 32'd58; 
32'd1971: dataIn2 = 32'd63; 
32'd1972: dataIn2 = 32'd78; 
32'd1973: dataIn2 = 32'd94; 
32'd1974: dataIn2 = 32'd50; 
32'd1975: dataIn2 = 32'd4; 
32'd1976: dataIn2 = 32'd27; 
32'd1977: dataIn2 = 32'd84; 
32'd1978: dataIn2 = 32'd79; 
32'd1979: dataIn2 = 32'd15; 
32'd1980: dataIn2 = 32'd33; 
32'd1981: dataIn2 = 32'd34; 
32'd1982: dataIn2 = 32'd84; 
32'd1983: dataIn2 = 32'd61; 
32'd1984: dataIn2 = 32'd60; 
32'd1985: dataIn2 = 32'd80; 
32'd1986: dataIn2 = 32'd9; 
32'd1987: dataIn2 = 32'd19; 
32'd1988: dataIn2 = 32'd53; 
32'd1989: dataIn2 = 32'd49; 
32'd1990: dataIn2 = 32'd89; 
32'd1991: dataIn2 = 32'd74; 
32'd1992: dataIn2 = 32'd7; 
32'd1993: dataIn2 = 32'd24; 
32'd1994: dataIn2 = 32'd65; 
32'd1995: dataIn2 = 32'd54; 
32'd1996: dataIn2 = 32'd61; 
32'd1997: dataIn2 = 32'd90; 
32'd1998: dataIn2 = 32'd50; 
32'd1999: dataIn2 = 32'd24; 
32'd2000: dataIn2 = 32'd34; 
32'd2001: dataIn2 = 32'd13; 
32'd2002: dataIn2 = 32'd88; 
32'd2003: dataIn2 = 32'd13; 
32'd2004: dataIn2 = 32'd70; 
32'd2005: dataIn2 = 32'd18; 
32'd2006: dataIn2 = 32'd18; 
32'd2007: dataIn2 = 32'd60; 
32'd2008: dataIn2 = 32'd17; 
32'd2009: dataIn2 = 32'd39; 
32'd2010: dataIn2 = 32'd38; 
32'd2011: dataIn2 = 32'd97; 
32'd2012: dataIn2 = 32'd95; 
32'd2013: dataIn2 = 32'd34; 
32'd2014: dataIn2 = 32'd98; 
32'd2015: dataIn2 = 32'd20; 
32'd2016: dataIn2 = 32'd43; 
32'd2017: dataIn2 = 32'd37; 
32'd2018: dataIn2 = 32'd73; 
32'd2019: dataIn2 = 32'd80; 
32'd2020: dataIn2 = 32'd63; 
32'd2021: dataIn2 = 32'd79; 
32'd2022: dataIn2 = 32'd68; 
32'd2023: dataIn2 = 32'd68; 
32'd2024: dataIn2 = 32'd63; 
32'd2025: dataIn2 = 32'd5; 
32'd2026: dataIn2 = 32'd1; 
32'd2027: dataIn2 = 32'd90; 
32'd2028: dataIn2 = 32'd88; 
32'd2029: dataIn2 = 32'd6; 
32'd2030: dataIn2 = 32'd55; 
32'd2031: dataIn2 = 32'd32; 
32'd2032: dataIn2 = 32'd49; 
32'd2033: dataIn2 = 32'd17; 
32'd2034: dataIn2 = 32'd29; 
32'd2035: dataIn2 = 32'd68; 
32'd2036: dataIn2 = 32'd81; 
32'd2037: dataIn2 = 32'd46; 
32'd2038: dataIn2 = 32'd18; 
32'd2039: dataIn2 = 32'd92; 
32'd2040: dataIn2 = 32'd23; 
32'd2041: dataIn2 = 32'd90; 
32'd2042: dataIn2 = 32'd32; 
32'd2043: dataIn2 = 32'd78; 
32'd2044: dataIn2 = 32'd9; 
32'd2045: dataIn2 = 32'd20; 
32'd2046: dataIn2 = 32'd79; 
32'd2047: dataIn2 = 32'd94; 
32'd2048: dataIn2 = 32'd37; 
32'd2049: dataIn2 = 32'd34; 
32'd2050: dataIn2 = 32'd25; 
32'd2051: dataIn2 = 32'd0; 
32'd2052: dataIn2 = 32'd38; 
32'd2053: dataIn2 = 32'd78; 
32'd2054: dataIn2 = 32'd74; 
32'd2055: dataIn2 = 32'd79; 
32'd2056: dataIn2 = 32'd98; 
32'd2057: dataIn2 = 32'd66; 
32'd2058: dataIn2 = 32'd65; 
32'd2059: dataIn2 = 32'd39; 
32'd2060: dataIn2 = 32'd43; 
32'd2061: dataIn2 = 32'd42; 
32'd2062: dataIn2 = 32'd61; 
32'd2063: dataIn2 = 32'd83; 
32'd2064: dataIn2 = 32'd96; 
32'd2065: dataIn2 = 32'd98; 
32'd2066: dataIn2 = 32'd27; 
32'd2067: dataIn2 = 32'd67; 
32'd2068: dataIn2 = 32'd82; 
32'd2069: dataIn2 = 32'd16; 
32'd2070: dataIn2 = 32'd6; 
32'd2071: dataIn2 = 32'd74; 
32'd2072: dataIn2 = 32'd63; 
32'd2073: dataIn2 = 32'd80; 
32'd2074: dataIn2 = 32'd87; 
32'd2075: dataIn2 = 32'd33; 
32'd2076: dataIn2 = 32'd11; 
32'd2077: dataIn2 = 32'd2; 
32'd2078: dataIn2 = 32'd74; 
32'd2079: dataIn2 = 32'd19; 
32'd2080: dataIn2 = 32'd78; 
32'd2081: dataIn2 = 32'd87; 
32'd2082: dataIn2 = 32'd1; 
32'd2083: dataIn2 = 32'd12; 
32'd2084: dataIn2 = 32'd41; 
32'd2085: dataIn2 = 32'd61; 
32'd2086: dataIn2 = 32'd9; 
32'd2087: dataIn2 = 32'd48; 
32'd2088: dataIn2 = 32'd85; 
32'd2089: dataIn2 = 32'd16; 
32'd2090: dataIn2 = 32'd52; 
32'd2091: dataIn2 = 32'd91; 
32'd2092: dataIn2 = 32'd15; 
32'd2093: dataIn2 = 32'd78; 
32'd2094: dataIn2 = 32'd85; 
32'd2095: dataIn2 = 32'd57; 
32'd2096: dataIn2 = 32'd73; 
32'd2097: dataIn2 = 32'd96; 
32'd2098: dataIn2 = 32'd44; 
32'd2099: dataIn2 = 32'd55; 
32'd2100: dataIn2 = 32'd65; 
32'd2101: dataIn2 = 32'd79; 
32'd2102: dataIn2 = 32'd62; 
32'd2103: dataIn2 = 32'd68; 
32'd2104: dataIn2 = 32'd12; 
32'd2105: dataIn2 = 32'd39; 
32'd2106: dataIn2 = 32'd94; 
32'd2107: dataIn2 = 32'd30; 
32'd2108: dataIn2 = 32'd64; 
32'd2109: dataIn2 = 32'd21; 
32'd2110: dataIn2 = 32'd0; 
32'd2111: dataIn2 = 32'd72; 
32'd2112: dataIn2 = 32'd44; 
32'd2113: dataIn2 = 32'd92; 
32'd2114: dataIn2 = 32'd95; 
32'd2115: dataIn2 = 32'd76; 
32'd2116: dataIn2 = 32'd46; 
32'd2117: dataIn2 = 32'd81; 
32'd2118: dataIn2 = 32'd28; 
32'd2119: dataIn2 = 32'd31; 
32'd2120: dataIn2 = 32'd79; 
32'd2121: dataIn2 = 32'd94; 
32'd2122: dataIn2 = 32'd95; 
32'd2123: dataIn2 = 32'd58; 
32'd2124: dataIn2 = 32'd11; 
32'd2125: dataIn2 = 32'd84; 
32'd2126: dataIn2 = 32'd69; 
32'd2127: dataIn2 = 32'd43; 
32'd2128: dataIn2 = 32'd5; 
32'd2129: dataIn2 = 32'd83; 
32'd2130: dataIn2 = 32'd26; 
32'd2131: dataIn2 = 32'd36; 
32'd2132: dataIn2 = 32'd71; 
32'd2133: dataIn2 = 32'd75; 
32'd2134: dataIn2 = 32'd4; 
32'd2135: dataIn2 = 32'd57; 
32'd2136: dataIn2 = 32'd43; 
32'd2137: dataIn2 = 32'd55; 
32'd2138: dataIn2 = 32'd14; 
32'd2139: dataIn2 = 32'd21; 
32'd2140: dataIn2 = 32'd13; 
32'd2141: dataIn2 = 32'd67; 
32'd2142: dataIn2 = 32'd61; 
32'd2143: dataIn2 = 32'd3; 
32'd2144: dataIn2 = 32'd48; 
32'd2145: dataIn2 = 32'd53; 
32'd2146: dataIn2 = 32'd42; 
32'd2147: dataIn2 = 32'd45; 
32'd2148: dataIn2 = 32'd89; 
32'd2149: dataIn2 = 32'd65; 
32'd2150: dataIn2 = 32'd38; 
32'd2151: dataIn2 = 32'd25; 
32'd2152: dataIn2 = 32'd92; 
32'd2153: dataIn2 = 32'd88; 
32'd2154: dataIn2 = 32'd47; 
32'd2155: dataIn2 = 32'd11; 
32'd2156: dataIn2 = 32'd3; 
32'd2157: dataIn2 = 32'd78; 
32'd2158: dataIn2 = 32'd80; 
32'd2159: dataIn2 = 32'd81; 
32'd2160: dataIn2 = 32'd55; 
32'd2161: dataIn2 = 32'd88; 
32'd2162: dataIn2 = 32'd96; 
32'd2163: dataIn2 = 32'd76; 
32'd2164: dataIn2 = 32'd46; 
32'd2165: dataIn2 = 32'd61; 
32'd2166: dataIn2 = 32'd12; 
32'd2167: dataIn2 = 32'd87; 
32'd2168: dataIn2 = 32'd50; 
32'd2169: dataIn2 = 32'd49; 
32'd2170: dataIn2 = 32'd55; 
32'd2171: dataIn2 = 32'd38; 
32'd2172: dataIn2 = 32'd32; 
32'd2173: dataIn2 = 32'd32; 
32'd2174: dataIn2 = 32'd51; 
32'd2175: dataIn2 = 32'd96; 
32'd2176: dataIn2 = 32'd7; 
32'd2177: dataIn2 = 32'd30; 
32'd2178: dataIn2 = 32'd16; 
32'd2179: dataIn2 = 32'd79; 
32'd2180: dataIn2 = 32'd35; 
32'd2181: dataIn2 = 32'd53; 
32'd2182: dataIn2 = 32'd51; 
32'd2183: dataIn2 = 32'd4; 
32'd2184: dataIn2 = 32'd11; 
32'd2185: dataIn2 = 32'd65; 
32'd2186: dataIn2 = 32'd44; 
32'd2187: dataIn2 = 32'd19; 
32'd2188: dataIn2 = 32'd100; 
32'd2189: dataIn2 = 32'd39; 
32'd2190: dataIn2 = 32'd34; 
32'd2191: dataIn2 = 32'd90; 
32'd2192: dataIn2 = 32'd34; 
32'd2193: dataIn2 = 32'd44; 
32'd2194: dataIn2 = 32'd49; 
32'd2195: dataIn2 = 32'd34; 
32'd2196: dataIn2 = 32'd70; 
32'd2197: dataIn2 = 32'd52; 
32'd2198: dataIn2 = 32'd50; 
32'd2199: dataIn2 = 32'd60; 
32'd2200: dataIn2 = 32'd84; 
32'd2201: dataIn2 = 32'd15; 
32'd2202: dataIn2 = 32'd87; 
32'd2203: dataIn2 = 32'd39; 
32'd2204: dataIn2 = 32'd81; 
32'd2205: dataIn2 = 32'd30; 
32'd2206: dataIn2 = 32'd60; 
32'd2207: dataIn2 = 32'd88; 
32'd2208: dataIn2 = 32'd27; 
32'd2209: dataIn2 = 32'd66; 
32'd2210: dataIn2 = 32'd96; 
32'd2211: dataIn2 = 32'd17; 
32'd2212: dataIn2 = 32'd22; 
32'd2213: dataIn2 = 32'd51; 
32'd2214: dataIn2 = 32'd47; 
32'd2215: dataIn2 = 32'd70; 
32'd2216: dataIn2 = 32'd19; 
32'd2217: dataIn2 = 32'd11; 
32'd2218: dataIn2 = 32'd83; 
32'd2219: dataIn2 = 32'd30; 
32'd2220: dataIn2 = 32'd95; 
32'd2221: dataIn2 = 32'd63; 
32'd2222: dataIn2 = 32'd82; 
32'd2223: dataIn2 = 32'd52; 
32'd2224: dataIn2 = 32'd73; 
32'd2225: dataIn2 = 32'd14; 
32'd2226: dataIn2 = 32'd16; 
32'd2227: dataIn2 = 32'd25; 
32'd2228: dataIn2 = 32'd61; 
32'd2229: dataIn2 = 32'd44; 
32'd2230: dataIn2 = 32'd83; 
32'd2231: dataIn2 = 32'd62; 
32'd2232: dataIn2 = 32'd42; 
32'd2233: dataIn2 = 32'd39; 
32'd2234: dataIn2 = 32'd14; 
32'd2235: dataIn2 = 32'd57; 
32'd2236: dataIn2 = 32'd17; 
32'd2237: dataIn2 = 32'd18; 
32'd2238: dataIn2 = 32'd90; 
32'd2239: dataIn2 = 32'd77; 
32'd2240: dataIn2 = 32'd24; 
32'd2241: dataIn2 = 32'd30; 
32'd2242: dataIn2 = 32'd75; 
32'd2243: dataIn2 = 32'd79; 
32'd2244: dataIn2 = 32'd17; 
32'd2245: dataIn2 = 32'd57; 
32'd2246: dataIn2 = 32'd51; 
32'd2247: dataIn2 = 32'd92; 
32'd2248: dataIn2 = 32'd1; 
32'd2249: dataIn2 = 32'd69; 
32'd2250: dataIn2 = 32'd2; 
32'd2251: dataIn2 = 32'd64; 
32'd2252: dataIn2 = 32'd99; 
32'd2253: dataIn2 = 32'd87; 
32'd2254: dataIn2 = 32'd93; 
32'd2255: dataIn2 = 32'd73; 
32'd2256: dataIn2 = 32'd30; 
32'd2257: dataIn2 = 32'd100; 
32'd2258: dataIn2 = 32'd44; 
32'd2259: dataIn2 = 32'd19; 
32'd2260: dataIn2 = 32'd42; 
32'd2261: dataIn2 = 32'd62; 
32'd2262: dataIn2 = 32'd90; 
32'd2263: dataIn2 = 32'd59; 
32'd2264: dataIn2 = 32'd45; 
32'd2265: dataIn2 = 32'd85; 
32'd2266: dataIn2 = 32'd48; 
32'd2267: dataIn2 = 32'd37; 
32'd2268: dataIn2 = 32'd35; 
32'd2269: dataIn2 = 32'd42; 
32'd2270: dataIn2 = 32'd56; 
32'd2271: dataIn2 = 32'd83; 
32'd2272: dataIn2 = 32'd94; 
32'd2273: dataIn2 = 32'd78; 
32'd2274: dataIn2 = 32'd20; 
32'd2275: dataIn2 = 32'd69; 
32'd2276: dataIn2 = 32'd14; 
32'd2277: dataIn2 = 32'd21; 
32'd2278: dataIn2 = 32'd70; 
32'd2279: dataIn2 = 32'd51; 
32'd2280: dataIn2 = 32'd2; 
32'd2281: dataIn2 = 32'd49; 
32'd2282: dataIn2 = 32'd6; 
32'd2283: dataIn2 = 32'd14; 
32'd2284: dataIn2 = 32'd20; 
32'd2285: dataIn2 = 32'd78; 
32'd2286: dataIn2 = 32'd78; 
32'd2287: dataIn2 = 32'd34; 
32'd2288: dataIn2 = 32'd59; 
32'd2289: dataIn2 = 32'd84; 
32'd2290: dataIn2 = 32'd77; 
32'd2291: dataIn2 = 32'd37; 
32'd2292: dataIn2 = 32'd0; 
32'd2293: dataIn2 = 32'd52; 
32'd2294: dataIn2 = 32'd22; 
32'd2295: dataIn2 = 32'd3; 
32'd2296: dataIn2 = 32'd48; 
32'd2297: dataIn2 = 32'd99; 
32'd2298: dataIn2 = 32'd94; 
32'd2299: dataIn2 = 32'd23; 
32'd2300: dataIn2 = 32'd50; 
32'd2301: dataIn2 = 32'd93; 
32'd2302: dataIn2 = 32'd89; 
32'd2303: dataIn2 = 32'd20; 
32'd2304: dataIn2 = 32'd20; 
32'd2305: dataIn2 = 32'd98; 
32'd2306: dataIn2 = 32'd38; 
32'd2307: dataIn2 = 32'd68; 
32'd2308: dataIn2 = 32'd17; 
32'd2309: dataIn2 = 32'd50; 
32'd2310: dataIn2 = 32'd64; 
32'd2311: dataIn2 = 32'd31; 
32'd2312: dataIn2 = 32'd44; 
32'd2313: dataIn2 = 32'd21; 
32'd2314: dataIn2 = 32'd42; 
32'd2315: dataIn2 = 32'd50; 
32'd2316: dataIn2 = 32'd40; 
32'd2317: dataIn2 = 32'd19; 
32'd2318: dataIn2 = 32'd59; 
32'd2319: dataIn2 = 32'd8; 
32'd2320: dataIn2 = 32'd74; 
32'd2321: dataIn2 = 32'd92; 
32'd2322: dataIn2 = 32'd20; 
32'd2323: dataIn2 = 32'd84; 
32'd2324: dataIn2 = 32'd82; 
32'd2325: dataIn2 = 32'd81; 
32'd2326: dataIn2 = 32'd2; 
32'd2327: dataIn2 = 32'd74; 
32'd2328: dataIn2 = 32'd51; 
32'd2329: dataIn2 = 32'd22; 
32'd2330: dataIn2 = 32'd68; 
32'd2331: dataIn2 = 32'd15; 
32'd2332: dataIn2 = 32'd43; 
32'd2333: dataIn2 = 32'd6; 
32'd2334: dataIn2 = 32'd5; 
32'd2335: dataIn2 = 32'd85; 
32'd2336: dataIn2 = 32'd89; 
32'd2337: dataIn2 = 32'd58; 
32'd2338: dataIn2 = 32'd89; 
32'd2339: dataIn2 = 32'd8; 
32'd2340: dataIn2 = 32'd32; 
32'd2341: dataIn2 = 32'd92; 
32'd2342: dataIn2 = 32'd89; 
32'd2343: dataIn2 = 32'd38; 
32'd2344: dataIn2 = 32'd65; 
32'd2345: dataIn2 = 32'd58; 
32'd2346: dataIn2 = 32'd41; 
32'd2347: dataIn2 = 32'd62; 
32'd2348: dataIn2 = 32'd87; 
32'd2349: dataIn2 = 32'd12; 
32'd2350: dataIn2 = 32'd44; 
32'd2351: dataIn2 = 32'd61; 
32'd2352: dataIn2 = 32'd79; 
32'd2353: dataIn2 = 32'd50; 
32'd2354: dataIn2 = 32'd61; 
32'd2355: dataIn2 = 32'd65; 
32'd2356: dataIn2 = 32'd45; 
32'd2357: dataIn2 = 32'd100; 
32'd2358: dataIn2 = 32'd13; 
32'd2359: dataIn2 = 32'd22; 
32'd2360: dataIn2 = 32'd80; 
32'd2361: dataIn2 = 32'd91; 
32'd2362: dataIn2 = 32'd0; 
32'd2363: dataIn2 = 32'd37; 
32'd2364: dataIn2 = 32'd100; 
32'd2365: dataIn2 = 32'd27; 
32'd2366: dataIn2 = 32'd26; 
32'd2367: dataIn2 = 32'd77; 
32'd2368: dataIn2 = 32'd89; 
32'd2369: dataIn2 = 32'd7; 
32'd2370: dataIn2 = 32'd81; 
32'd2371: dataIn2 = 32'd96; 
32'd2372: dataIn2 = 32'd79; 
32'd2373: dataIn2 = 32'd19; 
32'd2374: dataIn2 = 32'd61; 
32'd2375: dataIn2 = 32'd100; 
32'd2376: dataIn2 = 32'd35; 
32'd2377: dataIn2 = 32'd36; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_64_50.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
