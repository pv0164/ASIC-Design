//64x64 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 3277 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd330 ; 
  wdata_col_base = 32'd36070 ; 
  row_base = 32'd393470 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #343000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd393470: dataIn1 = 32'd0
; 
32'd393471: dataIn1 = 32'd50
; 
32'd393472: dataIn1 = 32'd100
; 
32'd393473: dataIn1 = 32'd150
; 
32'd393474: dataIn1 = 32'd193
; 
32'd393475: dataIn1 = 32'd243
; 
32'd393476: dataIn1 = 32'd294
; 
32'd393477: dataIn1 = 32'd347
; 
32'd393478: dataIn1 = 32'd394
; 
32'd393479: dataIn1 = 32'd441
; 
32'd393480: dataIn1 = 32'd489
; 
32'd393481: dataIn1 = 32'd539
; 
32'd393482: dataIn1 = 32'd588
; 
32'd393483: dataIn1 = 32'd639
; 
32'd393484: dataIn1 = 32'd692
; 
32'd393485: dataIn1 = 32'd742
; 
32'd393486: dataIn1 = 32'd790
; 
32'd393487: dataIn1 = 32'd835
; 
32'd393488: dataIn1 = 32'd887
; 
32'd393489: dataIn1 = 32'd939
; 
32'd393490: dataIn1 = 32'd992
; 
32'd393491: dataIn1 = 32'd1044
; 
32'd393492: dataIn1 = 32'd1097
; 
32'd393493: dataIn1 = 32'd1143
; 
32'd393494: dataIn1 = 32'd1189
; 
32'd393495: dataIn1 = 32'd1237
; 
32'd393496: dataIn1 = 32'd1283
; 
32'd393497: dataIn1 = 32'd1331
; 
32'd393498: dataIn1 = 32'd1377
; 
32'd393499: dataIn1 = 32'd1430
; 
32'd393500: dataIn1 = 32'd1481
; 
32'd393501: dataIn1 = 32'd1535
; 
32'd393502: dataIn1 = 32'd1585
; 
32'd393503: dataIn1 = 32'd1636
; 
32'd393504: dataIn1 = 32'd1683
; 
32'd393505: dataIn1 = 32'd1730
; 
32'd393506: dataIn1 = 32'd1784
; 
32'd393507: dataIn1 = 32'd1838
; 
32'd393508: dataIn1 = 32'd1885
; 
32'd393509: dataIn1 = 32'd1936
; 
32'd393510: dataIn1 = 32'd1984
; 
32'd393511: dataIn1 = 32'd2032
; 
32'd393512: dataIn1 = 32'd2086
; 
32'd393513: dataIn1 = 32'd2138
; 
32'd393514: dataIn1 = 32'd2187
; 
32'd393515: dataIn1 = 32'd2234
; 
32'd393516: dataIn1 = 32'd2280
; 
32'd393517: dataIn1 = 32'd2331
; 
32'd393518: dataIn1 = 32'd2384
; 
32'd393519: dataIn1 = 32'd2432
; 
32'd393520: dataIn1 = 32'd2480
; 
32'd393521: dataIn1 = 32'd2526
; 
32'd393522: dataIn1 = 32'd2574
; 
32'd393523: dataIn1 = 32'd2625
; 
32'd393524: dataIn1 = 32'd2676
; 
32'd393525: dataIn1 = 32'd2728
; 
32'd393526: dataIn1 = 32'd2779
; 
32'd393527: dataIn1 = 32'd2829
; 
32'd393528: dataIn1 = 32'd2877
; 
32'd393529: dataIn1 = 32'd2928
; 
32'd393530: dataIn1 = 32'd2979
; 
32'd393531: dataIn1 = 32'd3026
; 
32'd393532: dataIn1 = 32'd3076
; 
32'd393533: dataIn1 = 32'd3118
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd36070: dataIn1 = 32'd0
; 
32'd36071: dataIn1 = 32'd50
; 
32'd36072: dataIn1 = 32'd100
; 
32'd36073: dataIn1 = 32'd150
; 
32'd36074: dataIn1 = 32'd193
; 
32'd36075: dataIn1 = 32'd243
; 
32'd36076: dataIn1 = 32'd294
; 
32'd36077: dataIn1 = 32'd347
; 
32'd36078: dataIn1 = 32'd394
; 
32'd36079: dataIn1 = 32'd441
; 
32'd36080: dataIn1 = 32'd489
; 
32'd36081: dataIn1 = 32'd539
; 
32'd36082: dataIn1 = 32'd588
; 
32'd36083: dataIn1 = 32'd639
; 
32'd36084: dataIn1 = 32'd692
; 
32'd36085: dataIn1 = 32'd742
; 
32'd36086: dataIn1 = 32'd790
; 
32'd36087: dataIn1 = 32'd835
; 
32'd36088: dataIn1 = 32'd887
; 
32'd36089: dataIn1 = 32'd939
; 
32'd36090: dataIn1 = 32'd992
; 
32'd36091: dataIn1 = 32'd1044
; 
32'd36092: dataIn1 = 32'd1097
; 
32'd36093: dataIn1 = 32'd1143
; 
32'd36094: dataIn1 = 32'd1189
; 
32'd36095: dataIn1 = 32'd1237
; 
32'd36096: dataIn1 = 32'd1283
; 
32'd36097: dataIn1 = 32'd1331
; 
32'd36098: dataIn1 = 32'd1377
; 
32'd36099: dataIn1 = 32'd1430
; 
32'd36100: dataIn1 = 32'd1481
; 
32'd36101: dataIn1 = 32'd1535
; 
32'd36102: dataIn1 = 32'd1585
; 
32'd36103: dataIn1 = 32'd1636
; 
32'd36104: dataIn1 = 32'd1683
; 
32'd36105: dataIn1 = 32'd1730
; 
32'd36106: dataIn1 = 32'd1784
; 
32'd36107: dataIn1 = 32'd1838
; 
32'd36108: dataIn1 = 32'd1885
; 
32'd36109: dataIn1 = 32'd1936
; 
32'd36110: dataIn1 = 32'd1984
; 
32'd36111: dataIn1 = 32'd2032
; 
32'd36112: dataIn1 = 32'd2086
; 
32'd36113: dataIn1 = 32'd2138
; 
32'd36114: dataIn1 = 32'd2187
; 
32'd36115: dataIn1 = 32'd2234
; 
32'd36116: dataIn1 = 32'd2280
; 
32'd36117: dataIn1 = 32'd2331
; 
32'd36118: dataIn1 = 32'd2384
; 
32'd36119: dataIn1 = 32'd2432
; 
32'd36120: dataIn1 = 32'd2480
; 
32'd36121: dataIn1 = 32'd2526
; 
32'd36122: dataIn1 = 32'd2574
; 
32'd36123: dataIn1 = 32'd2625
; 
32'd36124: dataIn1 = 32'd2676
; 
32'd36125: dataIn1 = 32'd2728
; 
32'd36126: dataIn1 = 32'd2779
; 
32'd36127: dataIn1 = 32'd2829
; 
32'd36128: dataIn1 = 32'd2877
; 
32'd36129: dataIn1 = 32'd2928
; 
32'd36130: dataIn1 = 32'd2979
; 
32'd36131: dataIn1 = 32'd3026
; 
32'd36132: dataIn1 = 32'd3076
; 
32'd36133: dataIn1 = 32'd3118
; 
32'd36134: dataIn1 = 32'd3166
; 
32'd36135: dataIn1 = 32'd0
; 
32'd36136: dataIn1 = 32'd1
; 
32'd36137: dataIn1 = 32'd2
; 
32'd36138: dataIn1 = 32'd3
; 
32'd36139: dataIn1 = 32'd4
; 
32'd36140: dataIn1 = 32'd6
; 
32'd36141: dataIn1 = 32'd7
; 
32'd36142: dataIn1 = 32'd10
; 
32'd36143: dataIn1 = 32'd11
; 
32'd36144: dataIn1 = 32'd13
; 
32'd36145: dataIn1 = 32'd15
; 
32'd36146: dataIn1 = 32'd17
; 
32'd36147: dataIn1 = 32'd18
; 
32'd36148: dataIn1 = 32'd19
; 
32'd36149: dataIn1 = 32'd21
; 
32'd36150: dataIn1 = 32'd22
; 
32'd36151: dataIn1 = 32'd23
; 
32'd36152: dataIn1 = 32'd24
; 
32'd36153: dataIn1 = 32'd25
; 
32'd36154: dataIn1 = 32'd26
; 
32'd36155: dataIn1 = 32'd27
; 
32'd36156: dataIn1 = 32'd29
; 
32'd36157: dataIn1 = 32'd30
; 
32'd36158: dataIn1 = 32'd31
; 
32'd36159: dataIn1 = 32'd32
; 
32'd36160: dataIn1 = 32'd34
; 
32'd36161: dataIn1 = 32'd35
; 
32'd36162: dataIn1 = 32'd37
; 
32'd36163: dataIn1 = 32'd38
; 
32'd36164: dataIn1 = 32'd40
; 
32'd36165: dataIn1 = 32'd41
; 
32'd36166: dataIn1 = 32'd42
; 
32'd36167: dataIn1 = 32'd44
; 
32'd36168: dataIn1 = 32'd45
; 
32'd36169: dataIn1 = 32'd46
; 
32'd36170: dataIn1 = 32'd47
; 
32'd36171: dataIn1 = 32'd48
; 
32'd36172: dataIn1 = 32'd49
; 
32'd36173: dataIn1 = 32'd51
; 
32'd36174: dataIn1 = 32'd52
; 
32'd36175: dataIn1 = 32'd53
; 
32'd36176: dataIn1 = 32'd55
; 
32'd36177: dataIn1 = 32'd56
; 
32'd36178: dataIn1 = 32'd57
; 
32'd36179: dataIn1 = 32'd58
; 
32'd36180: dataIn1 = 32'd59
; 
32'd36181: dataIn1 = 32'd60
; 
32'd36182: dataIn1 = 32'd61
; 
32'd36183: dataIn1 = 32'd62
; 
32'd36184: dataIn1 = 32'd63
; 
32'd36185: dataIn1 = 32'd0
; 
32'd36186: dataIn1 = 32'd1
; 
32'd36187: dataIn1 = 32'd2
; 
32'd36188: dataIn1 = 32'd3
; 
32'd36189: dataIn1 = 32'd4
; 
32'd36190: dataIn1 = 32'd5
; 
32'd36191: dataIn1 = 32'd7
; 
32'd36192: dataIn1 = 32'd8
; 
32'd36193: dataIn1 = 32'd9
; 
32'd36194: dataIn1 = 32'd10
; 
32'd36195: dataIn1 = 32'd11
; 
32'd36196: dataIn1 = 32'd13
; 
32'd36197: dataIn1 = 32'd14
; 
32'd36198: dataIn1 = 32'd15
; 
32'd36199: dataIn1 = 32'd16
; 
32'd36200: dataIn1 = 32'd17
; 
32'd36201: dataIn1 = 32'd19
; 
32'd36202: dataIn1 = 32'd20
; 
32'd36203: dataIn1 = 32'd22
; 
32'd36204: dataIn1 = 32'd23
; 
32'd36205: dataIn1 = 32'd27
; 
32'd36206: dataIn1 = 32'd28
; 
32'd36207: dataIn1 = 32'd30
; 
32'd36208: dataIn1 = 32'd31
; 
32'd36209: dataIn1 = 32'd32
; 
32'd36210: dataIn1 = 32'd34
; 
32'd36211: dataIn1 = 32'd35
; 
32'd36212: dataIn1 = 32'd36
; 
32'd36213: dataIn1 = 32'd37
; 
32'd36214: dataIn1 = 32'd38
; 
32'd36215: dataIn1 = 32'd40
; 
32'd36216: dataIn1 = 32'd43
; 
32'd36217: dataIn1 = 32'd44
; 
32'd36218: dataIn1 = 32'd45
; 
32'd36219: dataIn1 = 32'd46
; 
32'd36220: dataIn1 = 32'd47
; 
32'd36221: dataIn1 = 32'd48
; 
32'd36222: dataIn1 = 32'd49
; 
32'd36223: dataIn1 = 32'd50
; 
32'd36224: dataIn1 = 32'd51
; 
32'd36225: dataIn1 = 32'd52
; 
32'd36226: dataIn1 = 32'd53
; 
32'd36227: dataIn1 = 32'd54
; 
32'd36228: dataIn1 = 32'd56
; 
32'd36229: dataIn1 = 32'd57
; 
32'd36230: dataIn1 = 32'd58
; 
32'd36231: dataIn1 = 32'd59
; 
32'd36232: dataIn1 = 32'd60
; 
32'd36233: dataIn1 = 32'd61
; 
32'd36234: dataIn1 = 32'd62
; 
32'd36235: dataIn1 = 32'd0
; 
32'd36236: dataIn1 = 32'd1
; 
32'd36237: dataIn1 = 32'd2
; 
32'd36238: dataIn1 = 32'd4
; 
32'd36239: dataIn1 = 32'd5
; 
32'd36240: dataIn1 = 32'd6
; 
32'd36241: dataIn1 = 32'd7
; 
32'd36242: dataIn1 = 32'd8
; 
32'd36243: dataIn1 = 32'd9
; 
32'd36244: dataIn1 = 32'd10
; 
32'd36245: dataIn1 = 32'd11
; 
32'd36246: dataIn1 = 32'd13
; 
32'd36247: dataIn1 = 32'd14
; 
32'd36248: dataIn1 = 32'd16
; 
32'd36249: dataIn1 = 32'd19
; 
32'd36250: dataIn1 = 32'd20
; 
32'd36251: dataIn1 = 32'd21
; 
32'd36252: dataIn1 = 32'd22
; 
32'd36253: dataIn1 = 32'd23
; 
32'd36254: dataIn1 = 32'd24
; 
32'd36255: dataIn1 = 32'd25
; 
32'd36256: dataIn1 = 32'd27
; 
32'd36257: dataIn1 = 32'd28
; 
32'd36258: dataIn1 = 32'd29
; 
32'd36259: dataIn1 = 32'd30
; 
32'd36260: dataIn1 = 32'd31
; 
32'd36261: dataIn1 = 32'd32
; 
32'd36262: dataIn1 = 32'd33
; 
32'd36263: dataIn1 = 32'd35
; 
32'd36264: dataIn1 = 32'd38
; 
32'd36265: dataIn1 = 32'd40
; 
32'd36266: dataIn1 = 32'd42
; 
32'd36267: dataIn1 = 32'd43
; 
32'd36268: dataIn1 = 32'd44
; 
32'd36269: dataIn1 = 32'd45
; 
32'd36270: dataIn1 = 32'd46
; 
32'd36271: dataIn1 = 32'd47
; 
32'd36272: dataIn1 = 32'd49
; 
32'd36273: dataIn1 = 32'd50
; 
32'd36274: dataIn1 = 32'd51
; 
32'd36275: dataIn1 = 32'd52
; 
32'd36276: dataIn1 = 32'd53
; 
32'd36277: dataIn1 = 32'd54
; 
32'd36278: dataIn1 = 32'd55
; 
32'd36279: dataIn1 = 32'd56
; 
32'd36280: dataIn1 = 32'd58
; 
32'd36281: dataIn1 = 32'd60
; 
32'd36282: dataIn1 = 32'd61
; 
32'd36283: dataIn1 = 32'd62
; 
32'd36284: dataIn1 = 32'd63
; 
32'd36285: dataIn1 = 32'd0
; 
32'd36286: dataIn1 = 32'd1
; 
32'd36287: dataIn1 = 32'd2
; 
32'd36288: dataIn1 = 32'd6
; 
32'd36289: dataIn1 = 32'd8
; 
32'd36290: dataIn1 = 32'd10
; 
32'd36291: dataIn1 = 32'd11
; 
32'd36292: dataIn1 = 32'd12
; 
32'd36293: dataIn1 = 32'd13
; 
32'd36294: dataIn1 = 32'd14
; 
32'd36295: dataIn1 = 32'd15
; 
32'd36296: dataIn1 = 32'd16
; 
32'd36297: dataIn1 = 32'd19
; 
32'd36298: dataIn1 = 32'd20
; 
32'd36299: dataIn1 = 32'd22
; 
32'd36300: dataIn1 = 32'd23
; 
32'd36301: dataIn1 = 32'd25
; 
32'd36302: dataIn1 = 32'd26
; 
32'd36303: dataIn1 = 32'd27
; 
32'd36304: dataIn1 = 32'd30
; 
32'd36305: dataIn1 = 32'd32
; 
32'd36306: dataIn1 = 32'd34
; 
32'd36307: dataIn1 = 32'd35
; 
32'd36308: dataIn1 = 32'd36
; 
32'd36309: dataIn1 = 32'd37
; 
32'd36310: dataIn1 = 32'd38
; 
32'd36311: dataIn1 = 32'd39
; 
32'd36312: dataIn1 = 32'd41
; 
32'd36313: dataIn1 = 32'd44
; 
32'd36314: dataIn1 = 32'd45
; 
32'd36315: dataIn1 = 32'd47
; 
32'd36316: dataIn1 = 32'd48
; 
32'd36317: dataIn1 = 32'd49
; 
32'd36318: dataIn1 = 32'd50
; 
32'd36319: dataIn1 = 32'd51
; 
32'd36320: dataIn1 = 32'd52
; 
32'd36321: dataIn1 = 32'd53
; 
32'd36322: dataIn1 = 32'd54
; 
32'd36323: dataIn1 = 32'd56
; 
32'd36324: dataIn1 = 32'd57
; 
32'd36325: dataIn1 = 32'd60
; 
32'd36326: dataIn1 = 32'd61
; 
32'd36327: dataIn1 = 32'd63
; 
32'd36328: dataIn1 = 32'd0
; 
32'd36329: dataIn1 = 32'd1
; 
32'd36330: dataIn1 = 32'd3
; 
32'd36331: dataIn1 = 32'd4
; 
32'd36332: dataIn1 = 32'd5
; 
32'd36333: dataIn1 = 32'd6
; 
32'd36334: dataIn1 = 32'd8
; 
32'd36335: dataIn1 = 32'd9
; 
32'd36336: dataIn1 = 32'd10
; 
32'd36337: dataIn1 = 32'd11
; 
32'd36338: dataIn1 = 32'd13
; 
32'd36339: dataIn1 = 32'd16
; 
32'd36340: dataIn1 = 32'd19
; 
32'd36341: dataIn1 = 32'd20
; 
32'd36342: dataIn1 = 32'd21
; 
32'd36343: dataIn1 = 32'd22
; 
32'd36344: dataIn1 = 32'd23
; 
32'd36345: dataIn1 = 32'd24
; 
32'd36346: dataIn1 = 32'd26
; 
32'd36347: dataIn1 = 32'd27
; 
32'd36348: dataIn1 = 32'd28
; 
32'd36349: dataIn1 = 32'd29
; 
32'd36350: dataIn1 = 32'd30
; 
32'd36351: dataIn1 = 32'd31
; 
32'd36352: dataIn1 = 32'd32
; 
32'd36353: dataIn1 = 32'd33
; 
32'd36354: dataIn1 = 32'd34
; 
32'd36355: dataIn1 = 32'd35
; 
32'd36356: dataIn1 = 32'd37
; 
32'd36357: dataIn1 = 32'd38
; 
32'd36358: dataIn1 = 32'd39
; 
32'd36359: dataIn1 = 32'd40
; 
32'd36360: dataIn1 = 32'd42
; 
32'd36361: dataIn1 = 32'd44
; 
32'd36362: dataIn1 = 32'd46
; 
32'd36363: dataIn1 = 32'd47
; 
32'd36364: dataIn1 = 32'd48
; 
32'd36365: dataIn1 = 32'd49
; 
32'd36366: dataIn1 = 32'd50
; 
32'd36367: dataIn1 = 32'd51
; 
32'd36368: dataIn1 = 32'd52
; 
32'd36369: dataIn1 = 32'd53
; 
32'd36370: dataIn1 = 32'd54
; 
32'd36371: dataIn1 = 32'd55
; 
32'd36372: dataIn1 = 32'd56
; 
32'd36373: dataIn1 = 32'd58
; 
32'd36374: dataIn1 = 32'd59
; 
32'd36375: dataIn1 = 32'd60
; 
32'd36376: dataIn1 = 32'd61
; 
32'd36377: dataIn1 = 32'd62
; 
32'd36378: dataIn1 = 32'd0
; 
32'd36379: dataIn1 = 32'd1
; 
32'd36380: dataIn1 = 32'd2
; 
32'd36381: dataIn1 = 32'd3
; 
32'd36382: dataIn1 = 32'd4
; 
32'd36383: dataIn1 = 32'd5
; 
32'd36384: dataIn1 = 32'd6
; 
32'd36385: dataIn1 = 32'd7
; 
32'd36386: dataIn1 = 32'd8
; 
32'd36387: dataIn1 = 32'd9
; 
32'd36388: dataIn1 = 32'd10
; 
32'd36389: dataIn1 = 32'd11
; 
32'd36390: dataIn1 = 32'd12
; 
32'd36391: dataIn1 = 32'd13
; 
32'd36392: dataIn1 = 32'd14
; 
32'd36393: dataIn1 = 32'd16
; 
32'd36394: dataIn1 = 32'd19
; 
32'd36395: dataIn1 = 32'd20
; 
32'd36396: dataIn1 = 32'd21
; 
32'd36397: dataIn1 = 32'd23
; 
32'd36398: dataIn1 = 32'd24
; 
32'd36399: dataIn1 = 32'd25
; 
32'd36400: dataIn1 = 32'd26
; 
32'd36401: dataIn1 = 32'd27
; 
32'd36402: dataIn1 = 32'd28
; 
32'd36403: dataIn1 = 32'd30
; 
32'd36404: dataIn1 = 32'd31
; 
32'd36405: dataIn1 = 32'd32
; 
32'd36406: dataIn1 = 32'd33
; 
32'd36407: dataIn1 = 32'd34
; 
32'd36408: dataIn1 = 32'd35
; 
32'd36409: dataIn1 = 32'd36
; 
32'd36410: dataIn1 = 32'd38
; 
32'd36411: dataIn1 = 32'd40
; 
32'd36412: dataIn1 = 32'd41
; 
32'd36413: dataIn1 = 32'd42
; 
32'd36414: dataIn1 = 32'd45
; 
32'd36415: dataIn1 = 32'd46
; 
32'd36416: dataIn1 = 32'd47
; 
32'd36417: dataIn1 = 32'd48
; 
32'd36418: dataIn1 = 32'd49
; 
32'd36419: dataIn1 = 32'd51
; 
32'd36420: dataIn1 = 32'd52
; 
32'd36421: dataIn1 = 32'd54
; 
32'd36422: dataIn1 = 32'd55
; 
32'd36423: dataIn1 = 32'd56
; 
32'd36424: dataIn1 = 32'd57
; 
32'd36425: dataIn1 = 32'd60
; 
32'd36426: dataIn1 = 32'd61
; 
32'd36427: dataIn1 = 32'd62
; 
32'd36428: dataIn1 = 32'd63
; 
32'd36429: dataIn1 = 32'd0
; 
32'd36430: dataIn1 = 32'd1
; 
32'd36431: dataIn1 = 32'd2
; 
32'd36432: dataIn1 = 32'd3
; 
32'd36433: dataIn1 = 32'd4
; 
32'd36434: dataIn1 = 32'd6
; 
32'd36435: dataIn1 = 32'd7
; 
32'd36436: dataIn1 = 32'd8
; 
32'd36437: dataIn1 = 32'd9
; 
32'd36438: dataIn1 = 32'd10
; 
32'd36439: dataIn1 = 32'd11
; 
32'd36440: dataIn1 = 32'd12
; 
32'd36441: dataIn1 = 32'd14
; 
32'd36442: dataIn1 = 32'd15
; 
32'd36443: dataIn1 = 32'd16
; 
32'd36444: dataIn1 = 32'd17
; 
32'd36445: dataIn1 = 32'd18
; 
32'd36446: dataIn1 = 32'd19
; 
32'd36447: dataIn1 = 32'd20
; 
32'd36448: dataIn1 = 32'd21
; 
32'd36449: dataIn1 = 32'd22
; 
32'd36450: dataIn1 = 32'd23
; 
32'd36451: dataIn1 = 32'd24
; 
32'd36452: dataIn1 = 32'd25
; 
32'd36453: dataIn1 = 32'd26
; 
32'd36454: dataIn1 = 32'd27
; 
32'd36455: dataIn1 = 32'd28
; 
32'd36456: dataIn1 = 32'd30
; 
32'd36457: dataIn1 = 32'd32
; 
32'd36458: dataIn1 = 32'd33
; 
32'd36459: dataIn1 = 32'd35
; 
32'd36460: dataIn1 = 32'd36
; 
32'd36461: dataIn1 = 32'd37
; 
32'd36462: dataIn1 = 32'd40
; 
32'd36463: dataIn1 = 32'd42
; 
32'd36464: dataIn1 = 32'd43
; 
32'd36465: dataIn1 = 32'd44
; 
32'd36466: dataIn1 = 32'd45
; 
32'd36467: dataIn1 = 32'd46
; 
32'd36468: dataIn1 = 32'd47
; 
32'd36469: dataIn1 = 32'd48
; 
32'd36470: dataIn1 = 32'd49
; 
32'd36471: dataIn1 = 32'd50
; 
32'd36472: dataIn1 = 32'd51
; 
32'd36473: dataIn1 = 32'd52
; 
32'd36474: dataIn1 = 32'd53
; 
32'd36475: dataIn1 = 32'd54
; 
32'd36476: dataIn1 = 32'd56
; 
32'd36477: dataIn1 = 32'd57
; 
32'd36478: dataIn1 = 32'd59
; 
32'd36479: dataIn1 = 32'd61
; 
32'd36480: dataIn1 = 32'd62
; 
32'd36481: dataIn1 = 32'd63
; 
32'd36482: dataIn1 = 32'd0
; 
32'd36483: dataIn1 = 32'd1
; 
32'd36484: dataIn1 = 32'd3
; 
32'd36485: dataIn1 = 32'd4
; 
32'd36486: dataIn1 = 32'd6
; 
32'd36487: dataIn1 = 32'd7
; 
32'd36488: dataIn1 = 32'd10
; 
32'd36489: dataIn1 = 32'd11
; 
32'd36490: dataIn1 = 32'd12
; 
32'd36491: dataIn1 = 32'd13
; 
32'd36492: dataIn1 = 32'd14
; 
32'd36493: dataIn1 = 32'd15
; 
32'd36494: dataIn1 = 32'd16
; 
32'd36495: dataIn1 = 32'd17
; 
32'd36496: dataIn1 = 32'd18
; 
32'd36497: dataIn1 = 32'd21
; 
32'd36498: dataIn1 = 32'd22
; 
32'd36499: dataIn1 = 32'd24
; 
32'd36500: dataIn1 = 32'd25
; 
32'd36501: dataIn1 = 32'd26
; 
32'd36502: dataIn1 = 32'd27
; 
32'd36503: dataIn1 = 32'd29
; 
32'd36504: dataIn1 = 32'd30
; 
32'd36505: dataIn1 = 32'd31
; 
32'd36506: dataIn1 = 32'd33
; 
32'd36507: dataIn1 = 32'd34
; 
32'd36508: dataIn1 = 32'd35
; 
32'd36509: dataIn1 = 32'd36
; 
32'd36510: dataIn1 = 32'd37
; 
32'd36511: dataIn1 = 32'd38
; 
32'd36512: dataIn1 = 32'd39
; 
32'd36513: dataIn1 = 32'd40
; 
32'd36514: dataIn1 = 32'd41
; 
32'd36515: dataIn1 = 32'd42
; 
32'd36516: dataIn1 = 32'd43
; 
32'd36517: dataIn1 = 32'd44
; 
32'd36518: dataIn1 = 32'd45
; 
32'd36519: dataIn1 = 32'd47
; 
32'd36520: dataIn1 = 32'd48
; 
32'd36521: dataIn1 = 32'd50
; 
32'd36522: dataIn1 = 32'd52
; 
32'd36523: dataIn1 = 32'd53
; 
32'd36524: dataIn1 = 32'd54
; 
32'd36525: dataIn1 = 32'd56
; 
32'd36526: dataIn1 = 32'd58
; 
32'd36527: dataIn1 = 32'd61
; 
32'd36528: dataIn1 = 32'd62
; 
32'd36529: dataIn1 = 32'd0
; 
32'd36530: dataIn1 = 32'd1
; 
32'd36531: dataIn1 = 32'd3
; 
32'd36532: dataIn1 = 32'd4
; 
32'd36533: dataIn1 = 32'd5
; 
32'd36534: dataIn1 = 32'd7
; 
32'd36535: dataIn1 = 32'd9
; 
32'd36536: dataIn1 = 32'd10
; 
32'd36537: dataIn1 = 32'd11
; 
32'd36538: dataIn1 = 32'd13
; 
32'd36539: dataIn1 = 32'd16
; 
32'd36540: dataIn1 = 32'd18
; 
32'd36541: dataIn1 = 32'd19
; 
32'd36542: dataIn1 = 32'd20
; 
32'd36543: dataIn1 = 32'd21
; 
32'd36544: dataIn1 = 32'd22
; 
32'd36545: dataIn1 = 32'd23
; 
32'd36546: dataIn1 = 32'd25
; 
32'd36547: dataIn1 = 32'd26
; 
32'd36548: dataIn1 = 32'd27
; 
32'd36549: dataIn1 = 32'd28
; 
32'd36550: dataIn1 = 32'd30
; 
32'd36551: dataIn1 = 32'd31
; 
32'd36552: dataIn1 = 32'd32
; 
32'd36553: dataIn1 = 32'd33
; 
32'd36554: dataIn1 = 32'd34
; 
32'd36555: dataIn1 = 32'd35
; 
32'd36556: dataIn1 = 32'd37
; 
32'd36557: dataIn1 = 32'd38
; 
32'd36558: dataIn1 = 32'd40
; 
32'd36559: dataIn1 = 32'd41
; 
32'd36560: dataIn1 = 32'd42
; 
32'd36561: dataIn1 = 32'd43
; 
32'd36562: dataIn1 = 32'd44
; 
32'd36563: dataIn1 = 32'd45
; 
32'd36564: dataIn1 = 32'd46
; 
32'd36565: dataIn1 = 32'd47
; 
32'd36566: dataIn1 = 32'd52
; 
32'd36567: dataIn1 = 32'd54
; 
32'd36568: dataIn1 = 32'd55
; 
32'd36569: dataIn1 = 32'd56
; 
32'd36570: dataIn1 = 32'd58
; 
32'd36571: dataIn1 = 32'd59
; 
32'd36572: dataIn1 = 32'd60
; 
32'd36573: dataIn1 = 32'd61
; 
32'd36574: dataIn1 = 32'd62
; 
32'd36575: dataIn1 = 32'd63
; 
32'd36576: dataIn1 = 32'd0
; 
32'd36577: dataIn1 = 32'd1
; 
32'd36578: dataIn1 = 32'd2
; 
32'd36579: dataIn1 = 32'd3
; 
32'd36580: dataIn1 = 32'd4
; 
32'd36581: dataIn1 = 32'd5
; 
32'd36582: dataIn1 = 32'd8
; 
32'd36583: dataIn1 = 32'd9
; 
32'd36584: dataIn1 = 32'd11
; 
32'd36585: dataIn1 = 32'd12
; 
32'd36586: dataIn1 = 32'd13
; 
32'd36587: dataIn1 = 32'd15
; 
32'd36588: dataIn1 = 32'd16
; 
32'd36589: dataIn1 = 32'd17
; 
32'd36590: dataIn1 = 32'd18
; 
32'd36591: dataIn1 = 32'd19
; 
32'd36592: dataIn1 = 32'd20
; 
32'd36593: dataIn1 = 32'd21
; 
32'd36594: dataIn1 = 32'd23
; 
32'd36595: dataIn1 = 32'd25
; 
32'd36596: dataIn1 = 32'd26
; 
32'd36597: dataIn1 = 32'd27
; 
32'd36598: dataIn1 = 32'd28
; 
32'd36599: dataIn1 = 32'd29
; 
32'd36600: dataIn1 = 32'd30
; 
32'd36601: dataIn1 = 32'd33
; 
32'd36602: dataIn1 = 32'd35
; 
32'd36603: dataIn1 = 32'd38
; 
32'd36604: dataIn1 = 32'd41
; 
32'd36605: dataIn1 = 32'd42
; 
32'd36606: dataIn1 = 32'd43
; 
32'd36607: dataIn1 = 32'd44
; 
32'd36608: dataIn1 = 32'd45
; 
32'd36609: dataIn1 = 32'd46
; 
32'd36610: dataIn1 = 32'd47
; 
32'd36611: dataIn1 = 32'd48
; 
32'd36612: dataIn1 = 32'd49
; 
32'd36613: dataIn1 = 32'd50
; 
32'd36614: dataIn1 = 32'd51
; 
32'd36615: dataIn1 = 32'd52
; 
32'd36616: dataIn1 = 32'd53
; 
32'd36617: dataIn1 = 32'd55
; 
32'd36618: dataIn1 = 32'd57
; 
32'd36619: dataIn1 = 32'd58
; 
32'd36620: dataIn1 = 32'd59
; 
32'd36621: dataIn1 = 32'd61
; 
32'd36622: dataIn1 = 32'd62
; 
32'd36623: dataIn1 = 32'd63
; 
32'd36624: dataIn1 = 32'd0
; 
32'd36625: dataIn1 = 32'd1
; 
32'd36626: dataIn1 = 32'd2
; 
32'd36627: dataIn1 = 32'd3
; 
32'd36628: dataIn1 = 32'd5
; 
32'd36629: dataIn1 = 32'd6
; 
32'd36630: dataIn1 = 32'd7
; 
32'd36631: dataIn1 = 32'd10
; 
32'd36632: dataIn1 = 32'd11
; 
32'd36633: dataIn1 = 32'd12
; 
32'd36634: dataIn1 = 32'd13
; 
32'd36635: dataIn1 = 32'd14
; 
32'd36636: dataIn1 = 32'd16
; 
32'd36637: dataIn1 = 32'd18
; 
32'd36638: dataIn1 = 32'd19
; 
32'd36639: dataIn1 = 32'd20
; 
32'd36640: dataIn1 = 32'd21
; 
32'd36641: dataIn1 = 32'd22
; 
32'd36642: dataIn1 = 32'd24
; 
32'd36643: dataIn1 = 32'd25
; 
32'd36644: dataIn1 = 32'd27
; 
32'd36645: dataIn1 = 32'd28
; 
32'd36646: dataIn1 = 32'd29
; 
32'd36647: dataIn1 = 32'd30
; 
32'd36648: dataIn1 = 32'd32
; 
32'd36649: dataIn1 = 32'd34
; 
32'd36650: dataIn1 = 32'd35
; 
32'd36651: dataIn1 = 32'd36
; 
32'd36652: dataIn1 = 32'd38
; 
32'd36653: dataIn1 = 32'd39
; 
32'd36654: dataIn1 = 32'd40
; 
32'd36655: dataIn1 = 32'd41
; 
32'd36656: dataIn1 = 32'd42
; 
32'd36657: dataIn1 = 32'd43
; 
32'd36658: dataIn1 = 32'd44
; 
32'd36659: dataIn1 = 32'd45
; 
32'd36660: dataIn1 = 32'd46
; 
32'd36661: dataIn1 = 32'd47
; 
32'd36662: dataIn1 = 32'd48
; 
32'd36663: dataIn1 = 32'd49
; 
32'd36664: dataIn1 = 32'd52
; 
32'd36665: dataIn1 = 32'd53
; 
32'd36666: dataIn1 = 32'd54
; 
32'd36667: dataIn1 = 32'd55
; 
32'd36668: dataIn1 = 32'd56
; 
32'd36669: dataIn1 = 32'd57
; 
32'd36670: dataIn1 = 32'd58
; 
32'd36671: dataIn1 = 32'd60
; 
32'd36672: dataIn1 = 32'd62
; 
32'd36673: dataIn1 = 32'd63
; 
32'd36674: dataIn1 = 32'd0
; 
32'd36675: dataIn1 = 32'd1
; 
32'd36676: dataIn1 = 32'd3
; 
32'd36677: dataIn1 = 32'd4
; 
32'd36678: dataIn1 = 32'd6
; 
32'd36679: dataIn1 = 32'd7
; 
32'd36680: dataIn1 = 32'd8
; 
32'd36681: dataIn1 = 32'd9
; 
32'd36682: dataIn1 = 32'd10
; 
32'd36683: dataIn1 = 32'd13
; 
32'd36684: dataIn1 = 32'd14
; 
32'd36685: dataIn1 = 32'd15
; 
32'd36686: dataIn1 = 32'd17
; 
32'd36687: dataIn1 = 32'd18
; 
32'd36688: dataIn1 = 32'd19
; 
32'd36689: dataIn1 = 32'd20
; 
32'd36690: dataIn1 = 32'd22
; 
32'd36691: dataIn1 = 32'd23
; 
32'd36692: dataIn1 = 32'd25
; 
32'd36693: dataIn1 = 32'd27
; 
32'd36694: dataIn1 = 32'd28
; 
32'd36695: dataIn1 = 32'd29
; 
32'd36696: dataIn1 = 32'd30
; 
32'd36697: dataIn1 = 32'd32
; 
32'd36698: dataIn1 = 32'd33
; 
32'd36699: dataIn1 = 32'd35
; 
32'd36700: dataIn1 = 32'd36
; 
32'd36701: dataIn1 = 32'd37
; 
32'd36702: dataIn1 = 32'd38
; 
32'd36703: dataIn1 = 32'd42
; 
32'd36704: dataIn1 = 32'd43
; 
32'd36705: dataIn1 = 32'd44
; 
32'd36706: dataIn1 = 32'd45
; 
32'd36707: dataIn1 = 32'd46
; 
32'd36708: dataIn1 = 32'd47
; 
32'd36709: dataIn1 = 32'd49
; 
32'd36710: dataIn1 = 32'd50
; 
32'd36711: dataIn1 = 32'd52
; 
32'd36712: dataIn1 = 32'd53
; 
32'd36713: dataIn1 = 32'd54
; 
32'd36714: dataIn1 = 32'd55
; 
32'd36715: dataIn1 = 32'd56
; 
32'd36716: dataIn1 = 32'd57
; 
32'd36717: dataIn1 = 32'd58
; 
32'd36718: dataIn1 = 32'd59
; 
32'd36719: dataIn1 = 32'd60
; 
32'd36720: dataIn1 = 32'd61
; 
32'd36721: dataIn1 = 32'd62
; 
32'd36722: dataIn1 = 32'd63
; 
32'd36723: dataIn1 = 32'd0
; 
32'd36724: dataIn1 = 32'd1
; 
32'd36725: dataIn1 = 32'd2
; 
32'd36726: dataIn1 = 32'd4
; 
32'd36727: dataIn1 = 32'd5
; 
32'd36728: dataIn1 = 32'd6
; 
32'd36729: dataIn1 = 32'd10
; 
32'd36730: dataIn1 = 32'd11
; 
32'd36731: dataIn1 = 32'd12
; 
32'd36732: dataIn1 = 32'd13
; 
32'd36733: dataIn1 = 32'd15
; 
32'd36734: dataIn1 = 32'd16
; 
32'd36735: dataIn1 = 32'd17
; 
32'd36736: dataIn1 = 32'd18
; 
32'd36737: dataIn1 = 32'd19
; 
32'd36738: dataIn1 = 32'd20
; 
32'd36739: dataIn1 = 32'd22
; 
32'd36740: dataIn1 = 32'd23
; 
32'd36741: dataIn1 = 32'd25
; 
32'd36742: dataIn1 = 32'd27
; 
32'd36743: dataIn1 = 32'd28
; 
32'd36744: dataIn1 = 32'd29
; 
32'd36745: dataIn1 = 32'd30
; 
32'd36746: dataIn1 = 32'd31
; 
32'd36747: dataIn1 = 32'd32
; 
32'd36748: dataIn1 = 32'd33
; 
32'd36749: dataIn1 = 32'd36
; 
32'd36750: dataIn1 = 32'd37
; 
32'd36751: dataIn1 = 32'd38
; 
32'd36752: dataIn1 = 32'd39
; 
32'd36753: dataIn1 = 32'd40
; 
32'd36754: dataIn1 = 32'd41
; 
32'd36755: dataIn1 = 32'd42
; 
32'd36756: dataIn1 = 32'd43
; 
32'd36757: dataIn1 = 32'd45
; 
32'd36758: dataIn1 = 32'd46
; 
32'd36759: dataIn1 = 32'd47
; 
32'd36760: dataIn1 = 32'd48
; 
32'd36761: dataIn1 = 32'd49
; 
32'd36762: dataIn1 = 32'd50
; 
32'd36763: dataIn1 = 32'd51
; 
32'd36764: dataIn1 = 32'd53
; 
32'd36765: dataIn1 = 32'd54
; 
32'd36766: dataIn1 = 32'd56
; 
32'd36767: dataIn1 = 32'd57
; 
32'd36768: dataIn1 = 32'd58
; 
32'd36769: dataIn1 = 32'd59
; 
32'd36770: dataIn1 = 32'd60
; 
32'd36771: dataIn1 = 32'd61
; 
32'd36772: dataIn1 = 32'd62
; 
32'd36773: dataIn1 = 32'd63
; 
32'd36774: dataIn1 = 32'd0
; 
32'd36775: dataIn1 = 32'd1
; 
32'd36776: dataIn1 = 32'd2
; 
32'd36777: dataIn1 = 32'd5
; 
32'd36778: dataIn1 = 32'd6
; 
32'd36779: dataIn1 = 32'd8
; 
32'd36780: dataIn1 = 32'd9
; 
32'd36781: dataIn1 = 32'd10
; 
32'd36782: dataIn1 = 32'd11
; 
32'd36783: dataIn1 = 32'd12
; 
32'd36784: dataIn1 = 32'd13
; 
32'd36785: dataIn1 = 32'd14
; 
32'd36786: dataIn1 = 32'd15
; 
32'd36787: dataIn1 = 32'd16
; 
32'd36788: dataIn1 = 32'd17
; 
32'd36789: dataIn1 = 32'd19
; 
32'd36790: dataIn1 = 32'd20
; 
32'd36791: dataIn1 = 32'd21
; 
32'd36792: dataIn1 = 32'd22
; 
32'd36793: dataIn1 = 32'd24
; 
32'd36794: dataIn1 = 32'd25
; 
32'd36795: dataIn1 = 32'd26
; 
32'd36796: dataIn1 = 32'd27
; 
32'd36797: dataIn1 = 32'd28
; 
32'd36798: dataIn1 = 32'd30
; 
32'd36799: dataIn1 = 32'd32
; 
32'd36800: dataIn1 = 32'd33
; 
32'd36801: dataIn1 = 32'd34
; 
32'd36802: dataIn1 = 32'd35
; 
32'd36803: dataIn1 = 32'd36
; 
32'd36804: dataIn1 = 32'd37
; 
32'd36805: dataIn1 = 32'd38
; 
32'd36806: dataIn1 = 32'd39
; 
32'd36807: dataIn1 = 32'd40
; 
32'd36808: dataIn1 = 32'd43
; 
32'd36809: dataIn1 = 32'd44
; 
32'd36810: dataIn1 = 32'd45
; 
32'd36811: dataIn1 = 32'd46
; 
32'd36812: dataIn1 = 32'd47
; 
32'd36813: dataIn1 = 32'd48
; 
32'd36814: dataIn1 = 32'd49
; 
32'd36815: dataIn1 = 32'd50
; 
32'd36816: dataIn1 = 32'd51
; 
32'd36817: dataIn1 = 32'd53
; 
32'd36818: dataIn1 = 32'd54
; 
32'd36819: dataIn1 = 32'd56
; 
32'd36820: dataIn1 = 32'd57
; 
32'd36821: dataIn1 = 32'd58
; 
32'd36822: dataIn1 = 32'd59
; 
32'd36823: dataIn1 = 32'd60
; 
32'd36824: dataIn1 = 32'd61
; 
32'd36825: dataIn1 = 32'd62
; 
32'd36826: dataIn1 = 32'd63
; 
32'd36827: dataIn1 = 32'd0
; 
32'd36828: dataIn1 = 32'd1
; 
32'd36829: dataIn1 = 32'd2
; 
32'd36830: dataIn1 = 32'd3
; 
32'd36831: dataIn1 = 32'd5
; 
32'd36832: dataIn1 = 32'd6
; 
32'd36833: dataIn1 = 32'd7
; 
32'd36834: dataIn1 = 32'd8
; 
32'd36835: dataIn1 = 32'd9
; 
32'd36836: dataIn1 = 32'd11
; 
32'd36837: dataIn1 = 32'd14
; 
32'd36838: dataIn1 = 32'd16
; 
32'd36839: dataIn1 = 32'd17
; 
32'd36840: dataIn1 = 32'd18
; 
32'd36841: dataIn1 = 32'd19
; 
32'd36842: dataIn1 = 32'd21
; 
32'd36843: dataIn1 = 32'd22
; 
32'd36844: dataIn1 = 32'd23
; 
32'd36845: dataIn1 = 32'd24
; 
32'd36846: dataIn1 = 32'd26
; 
32'd36847: dataIn1 = 32'd27
; 
32'd36848: dataIn1 = 32'd28
; 
32'd36849: dataIn1 = 32'd30
; 
32'd36850: dataIn1 = 32'd31
; 
32'd36851: dataIn1 = 32'd32
; 
32'd36852: dataIn1 = 32'd33
; 
32'd36853: dataIn1 = 32'd34
; 
32'd36854: dataIn1 = 32'd35
; 
32'd36855: dataIn1 = 32'd36
; 
32'd36856: dataIn1 = 32'd39
; 
32'd36857: dataIn1 = 32'd40
; 
32'd36858: dataIn1 = 32'd41
; 
32'd36859: dataIn1 = 32'd42
; 
32'd36860: dataIn1 = 32'd43
; 
32'd36861: dataIn1 = 32'd44
; 
32'd36862: dataIn1 = 32'd45
; 
32'd36863: dataIn1 = 32'd47
; 
32'd36864: dataIn1 = 32'd48
; 
32'd36865: dataIn1 = 32'd50
; 
32'd36866: dataIn1 = 32'd52
; 
32'd36867: dataIn1 = 32'd53
; 
32'd36868: dataIn1 = 32'd54
; 
32'd36869: dataIn1 = 32'd55
; 
32'd36870: dataIn1 = 32'd56
; 
32'd36871: dataIn1 = 32'd57
; 
32'd36872: dataIn1 = 32'd58
; 
32'd36873: dataIn1 = 32'd59
; 
32'd36874: dataIn1 = 32'd61
; 
32'd36875: dataIn1 = 32'd62
; 
32'd36876: dataIn1 = 32'd63
; 
32'd36877: dataIn1 = 32'd0
; 
32'd36878: dataIn1 = 32'd2
; 
32'd36879: dataIn1 = 32'd3
; 
32'd36880: dataIn1 = 32'd5
; 
32'd36881: dataIn1 = 32'd6
; 
32'd36882: dataIn1 = 32'd9
; 
32'd36883: dataIn1 = 32'd10
; 
32'd36884: dataIn1 = 32'd11
; 
32'd36885: dataIn1 = 32'd14
; 
32'd36886: dataIn1 = 32'd15
; 
32'd36887: dataIn1 = 32'd17
; 
32'd36888: dataIn1 = 32'd18
; 
32'd36889: dataIn1 = 32'd19
; 
32'd36890: dataIn1 = 32'd21
; 
32'd36891: dataIn1 = 32'd22
; 
32'd36892: dataIn1 = 32'd23
; 
32'd36893: dataIn1 = 32'd24
; 
32'd36894: dataIn1 = 32'd25
; 
32'd36895: dataIn1 = 32'd26
; 
32'd36896: dataIn1 = 32'd27
; 
32'd36897: dataIn1 = 32'd29
; 
32'd36898: dataIn1 = 32'd31
; 
32'd36899: dataIn1 = 32'd32
; 
32'd36900: dataIn1 = 32'd33
; 
32'd36901: dataIn1 = 32'd34
; 
32'd36902: dataIn1 = 32'd35
; 
32'd36903: dataIn1 = 32'd37
; 
32'd36904: dataIn1 = 32'd39
; 
32'd36905: dataIn1 = 32'd40
; 
32'd36906: dataIn1 = 32'd41
; 
32'd36907: dataIn1 = 32'd42
; 
32'd36908: dataIn1 = 32'd43
; 
32'd36909: dataIn1 = 32'd44
; 
32'd36910: dataIn1 = 32'd45
; 
32'd36911: dataIn1 = 32'd46
; 
32'd36912: dataIn1 = 32'd47
; 
32'd36913: dataIn1 = 32'd48
; 
32'd36914: dataIn1 = 32'd49
; 
32'd36915: dataIn1 = 32'd50
; 
32'd36916: dataIn1 = 32'd51
; 
32'd36917: dataIn1 = 32'd53
; 
32'd36918: dataIn1 = 32'd54
; 
32'd36919: dataIn1 = 32'd55
; 
32'd36920: dataIn1 = 32'd58
; 
32'd36921: dataIn1 = 32'd59
; 
32'd36922: dataIn1 = 32'd60
; 
32'd36923: dataIn1 = 32'd62
; 
32'd36924: dataIn1 = 32'd63
; 
32'd36925: dataIn1 = 32'd0
; 
32'd36926: dataIn1 = 32'd1
; 
32'd36927: dataIn1 = 32'd4
; 
32'd36928: dataIn1 = 32'd5
; 
32'd36929: dataIn1 = 32'd8
; 
32'd36930: dataIn1 = 32'd9
; 
32'd36931: dataIn1 = 32'd13
; 
32'd36932: dataIn1 = 32'd14
; 
32'd36933: dataIn1 = 32'd15
; 
32'd36934: dataIn1 = 32'd16
; 
32'd36935: dataIn1 = 32'd17
; 
32'd36936: dataIn1 = 32'd18
; 
32'd36937: dataIn1 = 32'd19
; 
32'd36938: dataIn1 = 32'd20
; 
32'd36939: dataIn1 = 32'd21
; 
32'd36940: dataIn1 = 32'd23
; 
32'd36941: dataIn1 = 32'd24
; 
32'd36942: dataIn1 = 32'd25
; 
32'd36943: dataIn1 = 32'd26
; 
32'd36944: dataIn1 = 32'd27
; 
32'd36945: dataIn1 = 32'd28
; 
32'd36946: dataIn1 = 32'd29
; 
32'd36947: dataIn1 = 32'd31
; 
32'd36948: dataIn1 = 32'd32
; 
32'd36949: dataIn1 = 32'd33
; 
32'd36950: dataIn1 = 32'd34
; 
32'd36951: dataIn1 = 32'd36
; 
32'd36952: dataIn1 = 32'd39
; 
32'd36953: dataIn1 = 32'd42
; 
32'd36954: dataIn1 = 32'd44
; 
32'd36955: dataIn1 = 32'd45
; 
32'd36956: dataIn1 = 32'd46
; 
32'd36957: dataIn1 = 32'd47
; 
32'd36958: dataIn1 = 32'd49
; 
32'd36959: dataIn1 = 32'd51
; 
32'd36960: dataIn1 = 32'd52
; 
32'd36961: dataIn1 = 32'd53
; 
32'd36962: dataIn1 = 32'd55
; 
32'd36963: dataIn1 = 32'd56
; 
32'd36964: dataIn1 = 32'd57
; 
32'd36965: dataIn1 = 32'd58
; 
32'd36966: dataIn1 = 32'd59
; 
32'd36967: dataIn1 = 32'd60
; 
32'd36968: dataIn1 = 32'd61
; 
32'd36969: dataIn1 = 32'd63
; 
32'd36970: dataIn1 = 32'd0
; 
32'd36971: dataIn1 = 32'd1
; 
32'd36972: dataIn1 = 32'd2
; 
32'd36973: dataIn1 = 32'd3
; 
32'd36974: dataIn1 = 32'd4
; 
32'd36975: dataIn1 = 32'd5
; 
32'd36976: dataIn1 = 32'd6
; 
32'd36977: dataIn1 = 32'd7
; 
32'd36978: dataIn1 = 32'd8
; 
32'd36979: dataIn1 = 32'd10
; 
32'd36980: dataIn1 = 32'd11
; 
32'd36981: dataIn1 = 32'd12
; 
32'd36982: dataIn1 = 32'd13
; 
32'd36983: dataIn1 = 32'd15
; 
32'd36984: dataIn1 = 32'd17
; 
32'd36985: dataIn1 = 32'd18
; 
32'd36986: dataIn1 = 32'd19
; 
32'd36987: dataIn1 = 32'd22
; 
32'd36988: dataIn1 = 32'd23
; 
32'd36989: dataIn1 = 32'd24
; 
32'd36990: dataIn1 = 32'd25
; 
32'd36991: dataIn1 = 32'd26
; 
32'd36992: dataIn1 = 32'd27
; 
32'd36993: dataIn1 = 32'd28
; 
32'd36994: dataIn1 = 32'd29
; 
32'd36995: dataIn1 = 32'd30
; 
32'd36996: dataIn1 = 32'd31
; 
32'd36997: dataIn1 = 32'd32
; 
32'd36998: dataIn1 = 32'd34
; 
32'd36999: dataIn1 = 32'd36
; 
32'd37000: dataIn1 = 32'd37
; 
32'd37001: dataIn1 = 32'd38
; 
32'd37002: dataIn1 = 32'd39
; 
32'd37003: dataIn1 = 32'd40
; 
32'd37004: dataIn1 = 32'd41
; 
32'd37005: dataIn1 = 32'd42
; 
32'd37006: dataIn1 = 32'd44
; 
32'd37007: dataIn1 = 32'd45
; 
32'd37008: dataIn1 = 32'd46
; 
32'd37009: dataIn1 = 32'd49
; 
32'd37010: dataIn1 = 32'd50
; 
32'd37011: dataIn1 = 32'd51
; 
32'd37012: dataIn1 = 32'd52
; 
32'd37013: dataIn1 = 32'd54
; 
32'd37014: dataIn1 = 32'd55
; 
32'd37015: dataIn1 = 32'd57
; 
32'd37016: dataIn1 = 32'd58
; 
32'd37017: dataIn1 = 32'd59
; 
32'd37018: dataIn1 = 32'd60
; 
32'd37019: dataIn1 = 32'd61
; 
32'd37020: dataIn1 = 32'd62
; 
32'd37021: dataIn1 = 32'd63
; 
32'd37022: dataIn1 = 32'd1
; 
32'd37023: dataIn1 = 32'd2
; 
32'd37024: dataIn1 = 32'd3
; 
32'd37025: dataIn1 = 32'd4
; 
32'd37026: dataIn1 = 32'd5
; 
32'd37027: dataIn1 = 32'd6
; 
32'd37028: dataIn1 = 32'd7
; 
32'd37029: dataIn1 = 32'd8
; 
32'd37030: dataIn1 = 32'd9
; 
32'd37031: dataIn1 = 32'd10
; 
32'd37032: dataIn1 = 32'd11
; 
32'd37033: dataIn1 = 32'd12
; 
32'd37034: dataIn1 = 32'd13
; 
32'd37035: dataIn1 = 32'd14
; 
32'd37036: dataIn1 = 32'd15
; 
32'd37037: dataIn1 = 32'd16
; 
32'd37038: dataIn1 = 32'd17
; 
32'd37039: dataIn1 = 32'd19
; 
32'd37040: dataIn1 = 32'd20
; 
32'd37041: dataIn1 = 32'd21
; 
32'd37042: dataIn1 = 32'd22
; 
32'd37043: dataIn1 = 32'd24
; 
32'd37044: dataIn1 = 32'd27
; 
32'd37045: dataIn1 = 32'd28
; 
32'd37046: dataIn1 = 32'd29
; 
32'd37047: dataIn1 = 32'd30
; 
32'd37048: dataIn1 = 32'd31
; 
32'd37049: dataIn1 = 32'd32
; 
32'd37050: dataIn1 = 32'd33
; 
32'd37051: dataIn1 = 32'd34
; 
32'd37052: dataIn1 = 32'd35
; 
32'd37053: dataIn1 = 32'd36
; 
32'd37054: dataIn1 = 32'd37
; 
32'd37055: dataIn1 = 32'd38
; 
32'd37056: dataIn1 = 32'd41
; 
32'd37057: dataIn1 = 32'd42
; 
32'd37058: dataIn1 = 32'd44
; 
32'd37059: dataIn1 = 32'd45
; 
32'd37060: dataIn1 = 32'd46
; 
32'd37061: dataIn1 = 32'd47
; 
32'd37062: dataIn1 = 32'd48
; 
32'd37063: dataIn1 = 32'd49
; 
32'd37064: dataIn1 = 32'd50
; 
32'd37065: dataIn1 = 32'd51
; 
32'd37066: dataIn1 = 32'd53
; 
32'd37067: dataIn1 = 32'd56
; 
32'd37068: dataIn1 = 32'd57
; 
32'd37069: dataIn1 = 32'd59
; 
32'd37070: dataIn1 = 32'd60
; 
32'd37071: dataIn1 = 32'd61
; 
32'd37072: dataIn1 = 32'd62
; 
32'd37073: dataIn1 = 32'd63
; 
32'd37074: dataIn1 = 32'd1
; 
32'd37075: dataIn1 = 32'd3
; 
32'd37076: dataIn1 = 32'd4
; 
32'd37077: dataIn1 = 32'd5
; 
32'd37078: dataIn1 = 32'd6
; 
32'd37079: dataIn1 = 32'd7
; 
32'd37080: dataIn1 = 32'd8
; 
32'd37081: dataIn1 = 32'd9
; 
32'd37082: dataIn1 = 32'd10
; 
32'd37083: dataIn1 = 32'd12
; 
32'd37084: dataIn1 = 32'd13
; 
32'd37085: dataIn1 = 32'd14
; 
32'd37086: dataIn1 = 32'd15
; 
32'd37087: dataIn1 = 32'd16
; 
32'd37088: dataIn1 = 32'd17
; 
32'd37089: dataIn1 = 32'd18
; 
32'd37090: dataIn1 = 32'd21
; 
32'd37091: dataIn1 = 32'd22
; 
32'd37092: dataIn1 = 32'd23
; 
32'd37093: dataIn1 = 32'd24
; 
32'd37094: dataIn1 = 32'd25
; 
32'd37095: dataIn1 = 32'd26
; 
32'd37096: dataIn1 = 32'd27
; 
32'd37097: dataIn1 = 32'd29
; 
32'd37098: dataIn1 = 32'd31
; 
32'd37099: dataIn1 = 32'd32
; 
32'd37100: dataIn1 = 32'd33
; 
32'd37101: dataIn1 = 32'd34
; 
32'd37102: dataIn1 = 32'd35
; 
32'd37103: dataIn1 = 32'd36
; 
32'd37104: dataIn1 = 32'd37
; 
32'd37105: dataIn1 = 32'd38
; 
32'd37106: dataIn1 = 32'd39
; 
32'd37107: dataIn1 = 32'd40
; 
32'd37108: dataIn1 = 32'd41
; 
32'd37109: dataIn1 = 32'd43
; 
32'd37110: dataIn1 = 32'd44
; 
32'd37111: dataIn1 = 32'd45
; 
32'd37112: dataIn1 = 32'd46
; 
32'd37113: dataIn1 = 32'd47
; 
32'd37114: dataIn1 = 32'd48
; 
32'd37115: dataIn1 = 32'd49
; 
32'd37116: dataIn1 = 32'd50
; 
32'd37117: dataIn1 = 32'd51
; 
32'd37118: dataIn1 = 32'd52
; 
32'd37119: dataIn1 = 32'd53
; 
32'd37120: dataIn1 = 32'd56
; 
32'd37121: dataIn1 = 32'd57
; 
32'd37122: dataIn1 = 32'd58
; 
32'd37123: dataIn1 = 32'd59
; 
32'd37124: dataIn1 = 32'd60
; 
32'd37125: dataIn1 = 32'd62
; 
32'd37126: dataIn1 = 32'd63
; 
32'd37127: dataIn1 = 32'd0
; 
32'd37128: dataIn1 = 32'd1
; 
32'd37129: dataIn1 = 32'd2
; 
32'd37130: dataIn1 = 32'd3
; 
32'd37131: dataIn1 = 32'd4
; 
32'd37132: dataIn1 = 32'd5
; 
32'd37133: dataIn1 = 32'd6
; 
32'd37134: dataIn1 = 32'd7
; 
32'd37135: dataIn1 = 32'd8
; 
32'd37136: dataIn1 = 32'd10
; 
32'd37137: dataIn1 = 32'd11
; 
32'd37138: dataIn1 = 32'd12
; 
32'd37139: dataIn1 = 32'd13
; 
32'd37140: dataIn1 = 32'd14
; 
32'd37141: dataIn1 = 32'd15
; 
32'd37142: dataIn1 = 32'd16
; 
32'd37143: dataIn1 = 32'd18
; 
32'd37144: dataIn1 = 32'd19
; 
32'd37145: dataIn1 = 32'd20
; 
32'd37146: dataIn1 = 32'd21
; 
32'd37147: dataIn1 = 32'd22
; 
32'd37148: dataIn1 = 32'd25
; 
32'd37149: dataIn1 = 32'd26
; 
32'd37150: dataIn1 = 32'd27
; 
32'd37151: dataIn1 = 32'd28
; 
32'd37152: dataIn1 = 32'd29
; 
32'd37153: dataIn1 = 32'd30
; 
32'd37154: dataIn1 = 32'd31
; 
32'd37155: dataIn1 = 32'd32
; 
32'd37156: dataIn1 = 32'd35
; 
32'd37157: dataIn1 = 32'd36
; 
32'd37158: dataIn1 = 32'd38
; 
32'd37159: dataIn1 = 32'd39
; 
32'd37160: dataIn1 = 32'd40
; 
32'd37161: dataIn1 = 32'd41
; 
32'd37162: dataIn1 = 32'd42
; 
32'd37163: dataIn1 = 32'd43
; 
32'd37164: dataIn1 = 32'd44
; 
32'd37165: dataIn1 = 32'd45
; 
32'd37166: dataIn1 = 32'd46
; 
32'd37167: dataIn1 = 32'd48
; 
32'd37168: dataIn1 = 32'd49
; 
32'd37169: dataIn1 = 32'd50
; 
32'd37170: dataIn1 = 32'd51
; 
32'd37171: dataIn1 = 32'd53
; 
32'd37172: dataIn1 = 32'd56
; 
32'd37173: dataIn1 = 32'd57
; 
32'd37174: dataIn1 = 32'd58
; 
32'd37175: dataIn1 = 32'd59
; 
32'd37176: dataIn1 = 32'd60
; 
32'd37177: dataIn1 = 32'd62
; 
32'd37178: dataIn1 = 32'd63
; 
32'd37179: dataIn1 = 32'd0
; 
32'd37180: dataIn1 = 32'd2
; 
32'd37181: dataIn1 = 32'd3
; 
32'd37182: dataIn1 = 32'd4
; 
32'd37183: dataIn1 = 32'd5
; 
32'd37184: dataIn1 = 32'd6
; 
32'd37185: dataIn1 = 32'd8
; 
32'd37186: dataIn1 = 32'd9
; 
32'd37187: dataIn1 = 32'd10
; 
32'd37188: dataIn1 = 32'd11
; 
32'd37189: dataIn1 = 32'd12
; 
32'd37190: dataIn1 = 32'd14
; 
32'd37191: dataIn1 = 32'd15
; 
32'd37192: dataIn1 = 32'd16
; 
32'd37193: dataIn1 = 32'd17
; 
32'd37194: dataIn1 = 32'd18
; 
32'd37195: dataIn1 = 32'd19
; 
32'd37196: dataIn1 = 32'd20
; 
32'd37197: dataIn1 = 32'd21
; 
32'd37198: dataIn1 = 32'd23
; 
32'd37199: dataIn1 = 32'd24
; 
32'd37200: dataIn1 = 32'd25
; 
32'd37201: dataIn1 = 32'd26
; 
32'd37202: dataIn1 = 32'd28
; 
32'd37203: dataIn1 = 32'd29
; 
32'd37204: dataIn1 = 32'd32
; 
32'd37205: dataIn1 = 32'd33
; 
32'd37206: dataIn1 = 32'd34
; 
32'd37207: dataIn1 = 32'd36
; 
32'd37208: dataIn1 = 32'd37
; 
32'd37209: dataIn1 = 32'd38
; 
32'd37210: dataIn1 = 32'd40
; 
32'd37211: dataIn1 = 32'd41
; 
32'd37212: dataIn1 = 32'd42
; 
32'd37213: dataIn1 = 32'd43
; 
32'd37214: dataIn1 = 32'd44
; 
32'd37215: dataIn1 = 32'd46
; 
32'd37216: dataIn1 = 32'd47
; 
32'd37217: dataIn1 = 32'd48
; 
32'd37218: dataIn1 = 32'd49
; 
32'd37219: dataIn1 = 32'd50
; 
32'd37220: dataIn1 = 32'd51
; 
32'd37221: dataIn1 = 32'd52
; 
32'd37222: dataIn1 = 32'd53
; 
32'd37223: dataIn1 = 32'd54
; 
32'd37224: dataIn1 = 32'd55
; 
32'd37225: dataIn1 = 32'd56
; 
32'd37226: dataIn1 = 32'd57
; 
32'd37227: dataIn1 = 32'd58
; 
32'd37228: dataIn1 = 32'd59
; 
32'd37229: dataIn1 = 32'd61
; 
32'd37230: dataIn1 = 32'd62
; 
32'd37231: dataIn1 = 32'd63
; 
32'd37232: dataIn1 = 32'd0
; 
32'd37233: dataIn1 = 32'd1
; 
32'd37234: dataIn1 = 32'd2
; 
32'd37235: dataIn1 = 32'd3
; 
32'd37236: dataIn1 = 32'd5
; 
32'd37237: dataIn1 = 32'd8
; 
32'd37238: dataIn1 = 32'd9
; 
32'd37239: dataIn1 = 32'd10
; 
32'd37240: dataIn1 = 32'd11
; 
32'd37241: dataIn1 = 32'd12
; 
32'd37242: dataIn1 = 32'd14
; 
32'd37243: dataIn1 = 32'd15
; 
32'd37244: dataIn1 = 32'd16
; 
32'd37245: dataIn1 = 32'd17
; 
32'd37246: dataIn1 = 32'd19
; 
32'd37247: dataIn1 = 32'd20
; 
32'd37248: dataIn1 = 32'd21
; 
32'd37249: dataIn1 = 32'd24
; 
32'd37250: dataIn1 = 32'd25
; 
32'd37251: dataIn1 = 32'd27
; 
32'd37252: dataIn1 = 32'd28
; 
32'd37253: dataIn1 = 32'd29
; 
32'd37254: dataIn1 = 32'd30
; 
32'd37255: dataIn1 = 32'd31
; 
32'd37256: dataIn1 = 32'd32
; 
32'd37257: dataIn1 = 32'd33
; 
32'd37258: dataIn1 = 32'd34
; 
32'd37259: dataIn1 = 32'd35
; 
32'd37260: dataIn1 = 32'd36
; 
32'd37261: dataIn1 = 32'd37
; 
32'd37262: dataIn1 = 32'd38
; 
32'd37263: dataIn1 = 32'd39
; 
32'd37264: dataIn1 = 32'd40
; 
32'd37265: dataIn1 = 32'd41
; 
32'd37266: dataIn1 = 32'd42
; 
32'd37267: dataIn1 = 32'd45
; 
32'd37268: dataIn1 = 32'd49
; 
32'd37269: dataIn1 = 32'd50
; 
32'd37270: dataIn1 = 32'd51
; 
32'd37271: dataIn1 = 32'd52
; 
32'd37272: dataIn1 = 32'd53
; 
32'd37273: dataIn1 = 32'd56
; 
32'd37274: dataIn1 = 32'd58
; 
32'd37275: dataIn1 = 32'd59
; 
32'd37276: dataIn1 = 32'd62
; 
32'd37277: dataIn1 = 32'd63
; 
32'd37278: dataIn1 = 32'd0
; 
32'd37279: dataIn1 = 32'd1
; 
32'd37280: dataIn1 = 32'd4
; 
32'd37281: dataIn1 = 32'd5
; 
32'd37282: dataIn1 = 32'd7
; 
32'd37283: dataIn1 = 32'd8
; 
32'd37284: dataIn1 = 32'd9
; 
32'd37285: dataIn1 = 32'd10
; 
32'd37286: dataIn1 = 32'd11
; 
32'd37287: dataIn1 = 32'd12
; 
32'd37288: dataIn1 = 32'd13
; 
32'd37289: dataIn1 = 32'd15
; 
32'd37290: dataIn1 = 32'd16
; 
32'd37291: dataIn1 = 32'd17
; 
32'd37292: dataIn1 = 32'd18
; 
32'd37293: dataIn1 = 32'd21
; 
32'd37294: dataIn1 = 32'd22
; 
32'd37295: dataIn1 = 32'd23
; 
32'd37296: dataIn1 = 32'd24
; 
32'd37297: dataIn1 = 32'd25
; 
32'd37298: dataIn1 = 32'd26
; 
32'd37299: dataIn1 = 32'd28
; 
32'd37300: dataIn1 = 32'd30
; 
32'd37301: dataIn1 = 32'd32
; 
32'd37302: dataIn1 = 32'd33
; 
32'd37303: dataIn1 = 32'd34
; 
32'd37304: dataIn1 = 32'd36
; 
32'd37305: dataIn1 = 32'd37
; 
32'd37306: dataIn1 = 32'd38
; 
32'd37307: dataIn1 = 32'd39
; 
32'd37308: dataIn1 = 32'd42
; 
32'd37309: dataIn1 = 32'd43
; 
32'd37310: dataIn1 = 32'd45
; 
32'd37311: dataIn1 = 32'd46
; 
32'd37312: dataIn1 = 32'd47
; 
32'd37313: dataIn1 = 32'd48
; 
32'd37314: dataIn1 = 32'd49
; 
32'd37315: dataIn1 = 32'd51
; 
32'd37316: dataIn1 = 32'd52
; 
32'd37317: dataIn1 = 32'd53
; 
32'd37318: dataIn1 = 32'd55
; 
32'd37319: dataIn1 = 32'd56
; 
32'd37320: dataIn1 = 32'd57
; 
32'd37321: dataIn1 = 32'd60
; 
32'd37322: dataIn1 = 32'd61
; 
32'd37323: dataIn1 = 32'd63
; 
32'd37324: dataIn1 = 32'd1
; 
32'd37325: dataIn1 = 32'd2
; 
32'd37326: dataIn1 = 32'd4
; 
32'd37327: dataIn1 = 32'd5
; 
32'd37328: dataIn1 = 32'd6
; 
32'd37329: dataIn1 = 32'd8
; 
32'd37330: dataIn1 = 32'd9
; 
32'd37331: dataIn1 = 32'd12
; 
32'd37332: dataIn1 = 32'd13
; 
32'd37333: dataIn1 = 32'd15
; 
32'd37334: dataIn1 = 32'd17
; 
32'd37335: dataIn1 = 32'd19
; 
32'd37336: dataIn1 = 32'd20
; 
32'd37337: dataIn1 = 32'd22
; 
32'd37338: dataIn1 = 32'd23
; 
32'd37339: dataIn1 = 32'd24
; 
32'd37340: dataIn1 = 32'd25
; 
32'd37341: dataIn1 = 32'd26
; 
32'd37342: dataIn1 = 32'd28
; 
32'd37343: dataIn1 = 32'd29
; 
32'd37344: dataIn1 = 32'd31
; 
32'd37345: dataIn1 = 32'd32
; 
32'd37346: dataIn1 = 32'd33
; 
32'd37347: dataIn1 = 32'd34
; 
32'd37348: dataIn1 = 32'd35
; 
32'd37349: dataIn1 = 32'd36
; 
32'd37350: dataIn1 = 32'd37
; 
32'd37351: dataIn1 = 32'd38
; 
32'd37352: dataIn1 = 32'd39
; 
32'd37353: dataIn1 = 32'd40
; 
32'd37354: dataIn1 = 32'd41
; 
32'd37355: dataIn1 = 32'd42
; 
32'd37356: dataIn1 = 32'd43
; 
32'd37357: dataIn1 = 32'd44
; 
32'd37358: dataIn1 = 32'd45
; 
32'd37359: dataIn1 = 32'd47
; 
32'd37360: dataIn1 = 32'd48
; 
32'd37361: dataIn1 = 32'd49
; 
32'd37362: dataIn1 = 32'd52
; 
32'd37363: dataIn1 = 32'd53
; 
32'd37364: dataIn1 = 32'd54
; 
32'd37365: dataIn1 = 32'd55
; 
32'd37366: dataIn1 = 32'd56
; 
32'd37367: dataIn1 = 32'd57
; 
32'd37368: dataIn1 = 32'd58
; 
32'd37369: dataIn1 = 32'd60
; 
32'd37370: dataIn1 = 32'd62
; 
32'd37371: dataIn1 = 32'd63
; 
32'd37372: dataIn1 = 32'd1
; 
32'd37373: dataIn1 = 32'd3
; 
32'd37374: dataIn1 = 32'd4
; 
32'd37375: dataIn1 = 32'd5
; 
32'd37376: dataIn1 = 32'd7
; 
32'd37377: dataIn1 = 32'd9
; 
32'd37378: dataIn1 = 32'd10
; 
32'd37379: dataIn1 = 32'd11
; 
32'd37380: dataIn1 = 32'd12
; 
32'd37381: dataIn1 = 32'd13
; 
32'd37382: dataIn1 = 32'd14
; 
32'd37383: dataIn1 = 32'd15
; 
32'd37384: dataIn1 = 32'd16
; 
32'd37385: dataIn1 = 32'd17
; 
32'd37386: dataIn1 = 32'd18
; 
32'd37387: dataIn1 = 32'd20
; 
32'd37388: dataIn1 = 32'd22
; 
32'd37389: dataIn1 = 32'd24
; 
32'd37390: dataIn1 = 32'd25
; 
32'd37391: dataIn1 = 32'd26
; 
32'd37392: dataIn1 = 32'd27
; 
32'd37393: dataIn1 = 32'd28
; 
32'd37394: dataIn1 = 32'd29
; 
32'd37395: dataIn1 = 32'd30
; 
32'd37396: dataIn1 = 32'd33
; 
32'd37397: dataIn1 = 32'd34
; 
32'd37398: dataIn1 = 32'd35
; 
32'd37399: dataIn1 = 32'd36
; 
32'd37400: dataIn1 = 32'd37
; 
32'd37401: dataIn1 = 32'd38
; 
32'd37402: dataIn1 = 32'd39
; 
32'd37403: dataIn1 = 32'd41
; 
32'd37404: dataIn1 = 32'd42
; 
32'd37405: dataIn1 = 32'd45
; 
32'd37406: dataIn1 = 32'd46
; 
32'd37407: dataIn1 = 32'd48
; 
32'd37408: dataIn1 = 32'd49
; 
32'd37409: dataIn1 = 32'd50
; 
32'd37410: dataIn1 = 32'd53
; 
32'd37411: dataIn1 = 32'd55
; 
32'd37412: dataIn1 = 32'd56
; 
32'd37413: dataIn1 = 32'd57
; 
32'd37414: dataIn1 = 32'd58
; 
32'd37415: dataIn1 = 32'd59
; 
32'd37416: dataIn1 = 32'd60
; 
32'd37417: dataIn1 = 32'd62
; 
32'd37418: dataIn1 = 32'd0
; 
32'd37419: dataIn1 = 32'd1
; 
32'd37420: dataIn1 = 32'd2
; 
32'd37421: dataIn1 = 32'd3
; 
32'd37422: dataIn1 = 32'd4
; 
32'd37423: dataIn1 = 32'd5
; 
32'd37424: dataIn1 = 32'd8
; 
32'd37425: dataIn1 = 32'd9
; 
32'd37426: dataIn1 = 32'd10
; 
32'd37427: dataIn1 = 32'd11
; 
32'd37428: dataIn1 = 32'd12
; 
32'd37429: dataIn1 = 32'd13
; 
32'd37430: dataIn1 = 32'd17
; 
32'd37431: dataIn1 = 32'd18
; 
32'd37432: dataIn1 = 32'd19
; 
32'd37433: dataIn1 = 32'd20
; 
32'd37434: dataIn1 = 32'd21
; 
32'd37435: dataIn1 = 32'd22
; 
32'd37436: dataIn1 = 32'd24
; 
32'd37437: dataIn1 = 32'd25
; 
32'd37438: dataIn1 = 32'd26
; 
32'd37439: dataIn1 = 32'd27
; 
32'd37440: dataIn1 = 32'd28
; 
32'd37441: dataIn1 = 32'd29
; 
32'd37442: dataIn1 = 32'd30
; 
32'd37443: dataIn1 = 32'd31
; 
32'd37444: dataIn1 = 32'd32
; 
32'd37445: dataIn1 = 32'd35
; 
32'd37446: dataIn1 = 32'd37
; 
32'd37447: dataIn1 = 32'd38
; 
32'd37448: dataIn1 = 32'd39
; 
32'd37449: dataIn1 = 32'd40
; 
32'd37450: dataIn1 = 32'd41
; 
32'd37451: dataIn1 = 32'd42
; 
32'd37452: dataIn1 = 32'd44
; 
32'd37453: dataIn1 = 32'd45
; 
32'd37454: dataIn1 = 32'd46
; 
32'd37455: dataIn1 = 32'd49
; 
32'd37456: dataIn1 = 32'd50
; 
32'd37457: dataIn1 = 32'd51
; 
32'd37458: dataIn1 = 32'd52
; 
32'd37459: dataIn1 = 32'd53
; 
32'd37460: dataIn1 = 32'd54
; 
32'd37461: dataIn1 = 32'd57
; 
32'd37462: dataIn1 = 32'd58
; 
32'd37463: dataIn1 = 32'd60
; 
32'd37464: dataIn1 = 32'd61
; 
32'd37465: dataIn1 = 32'd62
; 
32'd37466: dataIn1 = 32'd1
; 
32'd37467: dataIn1 = 32'd2
; 
32'd37468: dataIn1 = 32'd3
; 
32'd37469: dataIn1 = 32'd5
; 
32'd37470: dataIn1 = 32'd7
; 
32'd37471: dataIn1 = 32'd8
; 
32'd37472: dataIn1 = 32'd9
; 
32'd37473: dataIn1 = 32'd10
; 
32'd37474: dataIn1 = 32'd13
; 
32'd37475: dataIn1 = 32'd16
; 
32'd37476: dataIn1 = 32'd17
; 
32'd37477: dataIn1 = 32'd18
; 
32'd37478: dataIn1 = 32'd20
; 
32'd37479: dataIn1 = 32'd21
; 
32'd37480: dataIn1 = 32'd24
; 
32'd37481: dataIn1 = 32'd25
; 
32'd37482: dataIn1 = 32'd26
; 
32'd37483: dataIn1 = 32'd27
; 
32'd37484: dataIn1 = 32'd28
; 
32'd37485: dataIn1 = 32'd30
; 
32'd37486: dataIn1 = 32'd31
; 
32'd37487: dataIn1 = 32'd32
; 
32'd37488: dataIn1 = 32'd33
; 
32'd37489: dataIn1 = 32'd34
; 
32'd37490: dataIn1 = 32'd35
; 
32'd37491: dataIn1 = 32'd36
; 
32'd37492: dataIn1 = 32'd38
; 
32'd37493: dataIn1 = 32'd39
; 
32'd37494: dataIn1 = 32'd40
; 
32'd37495: dataIn1 = 32'd43
; 
32'd37496: dataIn1 = 32'd44
; 
32'd37497: dataIn1 = 32'd45
; 
32'd37498: dataIn1 = 32'd46
; 
32'd37499: dataIn1 = 32'd47
; 
32'd37500: dataIn1 = 32'd48
; 
32'd37501: dataIn1 = 32'd51
; 
32'd37502: dataIn1 = 32'd52
; 
32'd37503: dataIn1 = 32'd54
; 
32'd37504: dataIn1 = 32'd55
; 
32'd37505: dataIn1 = 32'd56
; 
32'd37506: dataIn1 = 32'd58
; 
32'd37507: dataIn1 = 32'd59
; 
32'd37508: dataIn1 = 32'd60
; 
32'd37509: dataIn1 = 32'd61
; 
32'd37510: dataIn1 = 32'd62
; 
32'd37511: dataIn1 = 32'd63
; 
32'd37512: dataIn1 = 32'd0
; 
32'd37513: dataIn1 = 32'd1
; 
32'd37514: dataIn1 = 32'd2
; 
32'd37515: dataIn1 = 32'd3
; 
32'd37516: dataIn1 = 32'd4
; 
32'd37517: dataIn1 = 32'd5
; 
32'd37518: dataIn1 = 32'd6
; 
32'd37519: dataIn1 = 32'd7
; 
32'd37520: dataIn1 = 32'd8
; 
32'd37521: dataIn1 = 32'd10
; 
32'd37522: dataIn1 = 32'd11
; 
32'd37523: dataIn1 = 32'd12
; 
32'd37524: dataIn1 = 32'd14
; 
32'd37525: dataIn1 = 32'd15
; 
32'd37526: dataIn1 = 32'd17
; 
32'd37527: dataIn1 = 32'd18
; 
32'd37528: dataIn1 = 32'd19
; 
32'd37529: dataIn1 = 32'd21
; 
32'd37530: dataIn1 = 32'd22
; 
32'd37531: dataIn1 = 32'd23
; 
32'd37532: dataIn1 = 32'd24
; 
32'd37533: dataIn1 = 32'd25
; 
32'd37534: dataIn1 = 32'd26
; 
32'd37535: dataIn1 = 32'd27
; 
32'd37536: dataIn1 = 32'd28
; 
32'd37537: dataIn1 = 32'd30
; 
32'd37538: dataIn1 = 32'd31
; 
32'd37539: dataIn1 = 32'd32
; 
32'd37540: dataIn1 = 32'd33
; 
32'd37541: dataIn1 = 32'd34
; 
32'd37542: dataIn1 = 32'd35
; 
32'd37543: dataIn1 = 32'd38
; 
32'd37544: dataIn1 = 32'd39
; 
32'd37545: dataIn1 = 32'd40
; 
32'd37546: dataIn1 = 32'd41
; 
32'd37547: dataIn1 = 32'd42
; 
32'd37548: dataIn1 = 32'd43
; 
32'd37549: dataIn1 = 32'd44
; 
32'd37550: dataIn1 = 32'd46
; 
32'd37551: dataIn1 = 32'd47
; 
32'd37552: dataIn1 = 32'd49
; 
32'd37553: dataIn1 = 32'd50
; 
32'd37554: dataIn1 = 32'd51
; 
32'd37555: dataIn1 = 32'd52
; 
32'd37556: dataIn1 = 32'd53
; 
32'd37557: dataIn1 = 32'd54
; 
32'd37558: dataIn1 = 32'd56
; 
32'd37559: dataIn1 = 32'd57
; 
32'd37560: dataIn1 = 32'd58
; 
32'd37561: dataIn1 = 32'd59
; 
32'd37562: dataIn1 = 32'd60
; 
32'd37563: dataIn1 = 32'd61
; 
32'd37564: dataIn1 = 32'd62
; 
32'd37565: dataIn1 = 32'd0
; 
32'd37566: dataIn1 = 32'd1
; 
32'd37567: dataIn1 = 32'd3
; 
32'd37568: dataIn1 = 32'd4
; 
32'd37569: dataIn1 = 32'd5
; 
32'd37570: dataIn1 = 32'd7
; 
32'd37571: dataIn1 = 32'd9
; 
32'd37572: dataIn1 = 32'd10
; 
32'd37573: dataIn1 = 32'd11
; 
32'd37574: dataIn1 = 32'd13
; 
32'd37575: dataIn1 = 32'd15
; 
32'd37576: dataIn1 = 32'd16
; 
32'd37577: dataIn1 = 32'd17
; 
32'd37578: dataIn1 = 32'd18
; 
32'd37579: dataIn1 = 32'd19
; 
32'd37580: dataIn1 = 32'd20
; 
32'd37581: dataIn1 = 32'd21
; 
32'd37582: dataIn1 = 32'd22
; 
32'd37583: dataIn1 = 32'd23
; 
32'd37584: dataIn1 = 32'd25
; 
32'd37585: dataIn1 = 32'd26
; 
32'd37586: dataIn1 = 32'd27
; 
32'd37587: dataIn1 = 32'd28
; 
32'd37588: dataIn1 = 32'd29
; 
32'd37589: dataIn1 = 32'd30
; 
32'd37590: dataIn1 = 32'd31
; 
32'd37591: dataIn1 = 32'd32
; 
32'd37592: dataIn1 = 32'd34
; 
32'd37593: dataIn1 = 32'd36
; 
32'd37594: dataIn1 = 32'd37
; 
32'd37595: dataIn1 = 32'd39
; 
32'd37596: dataIn1 = 32'd40
; 
32'd37597: dataIn1 = 32'd41
; 
32'd37598: dataIn1 = 32'd42
; 
32'd37599: dataIn1 = 32'd44
; 
32'd37600: dataIn1 = 32'd45
; 
32'd37601: dataIn1 = 32'd47
; 
32'd37602: dataIn1 = 32'd48
; 
32'd37603: dataIn1 = 32'd49
; 
32'd37604: dataIn1 = 32'd50
; 
32'd37605: dataIn1 = 32'd51
; 
32'd37606: dataIn1 = 32'd52
; 
32'd37607: dataIn1 = 32'd53
; 
32'd37608: dataIn1 = 32'd54
; 
32'd37609: dataIn1 = 32'd55
; 
32'd37610: dataIn1 = 32'd56
; 
32'd37611: dataIn1 = 32'd58
; 
32'd37612: dataIn1 = 32'd60
; 
32'd37613: dataIn1 = 32'd61
; 
32'd37614: dataIn1 = 32'd62
; 
32'd37615: dataIn1 = 32'd63
; 
32'd37616: dataIn1 = 32'd0
; 
32'd37617: dataIn1 = 32'd1
; 
32'd37618: dataIn1 = 32'd2
; 
32'd37619: dataIn1 = 32'd3
; 
32'd37620: dataIn1 = 32'd4
; 
32'd37621: dataIn1 = 32'd5
; 
32'd37622: dataIn1 = 32'd6
; 
32'd37623: dataIn1 = 32'd7
; 
32'd37624: dataIn1 = 32'd8
; 
32'd37625: dataIn1 = 32'd10
; 
32'd37626: dataIn1 = 32'd12
; 
32'd37627: dataIn1 = 32'd13
; 
32'd37628: dataIn1 = 32'd14
; 
32'd37629: dataIn1 = 32'd15
; 
32'd37630: dataIn1 = 32'd16
; 
32'd37631: dataIn1 = 32'd18
; 
32'd37632: dataIn1 = 32'd21
; 
32'd37633: dataIn1 = 32'd22
; 
32'd37634: dataIn1 = 32'd23
; 
32'd37635: dataIn1 = 32'd24
; 
32'd37636: dataIn1 = 32'd27
; 
32'd37637: dataIn1 = 32'd29
; 
32'd37638: dataIn1 = 32'd30
; 
32'd37639: dataIn1 = 32'd31
; 
32'd37640: dataIn1 = 32'd32
; 
32'd37641: dataIn1 = 32'd33
; 
32'd37642: dataIn1 = 32'd34
; 
32'd37643: dataIn1 = 32'd35
; 
32'd37644: dataIn1 = 32'd36
; 
32'd37645: dataIn1 = 32'd37
; 
32'd37646: dataIn1 = 32'd39
; 
32'd37647: dataIn1 = 32'd40
; 
32'd37648: dataIn1 = 32'd41
; 
32'd37649: dataIn1 = 32'd42
; 
32'd37650: dataIn1 = 32'd43
; 
32'd37651: dataIn1 = 32'd44
; 
32'd37652: dataIn1 = 32'd45
; 
32'd37653: dataIn1 = 32'd46
; 
32'd37654: dataIn1 = 32'd48
; 
32'd37655: dataIn1 = 32'd49
; 
32'd37656: dataIn1 = 32'd50
; 
32'd37657: dataIn1 = 32'd51
; 
32'd37658: dataIn1 = 32'd52
; 
32'd37659: dataIn1 = 32'd53
; 
32'd37660: dataIn1 = 32'd54
; 
32'd37661: dataIn1 = 32'd55
; 
32'd37662: dataIn1 = 32'd56
; 
32'd37663: dataIn1 = 32'd57
; 
32'd37664: dataIn1 = 32'd58
; 
32'd37665: dataIn1 = 32'd59
; 
32'd37666: dataIn1 = 32'd60
; 
32'd37667: dataIn1 = 32'd61
; 
32'd37668: dataIn1 = 32'd62
; 
32'd37669: dataIn1 = 32'd63
; 
32'd37670: dataIn1 = 32'd0
; 
32'd37671: dataIn1 = 32'd1
; 
32'd37672: dataIn1 = 32'd3
; 
32'd37673: dataIn1 = 32'd5
; 
32'd37674: dataIn1 = 32'd7
; 
32'd37675: dataIn1 = 32'd9
; 
32'd37676: dataIn1 = 32'd10
; 
32'd37677: dataIn1 = 32'd11
; 
32'd37678: dataIn1 = 32'd12
; 
32'd37679: dataIn1 = 32'd13
; 
32'd37680: dataIn1 = 32'd14
; 
32'd37681: dataIn1 = 32'd15
; 
32'd37682: dataIn1 = 32'd17
; 
32'd37683: dataIn1 = 32'd18
; 
32'd37684: dataIn1 = 32'd20
; 
32'd37685: dataIn1 = 32'd22
; 
32'd37686: dataIn1 = 32'd23
; 
32'd37687: dataIn1 = 32'd24
; 
32'd37688: dataIn1 = 32'd26
; 
32'd37689: dataIn1 = 32'd28
; 
32'd37690: dataIn1 = 32'd29
; 
32'd37691: dataIn1 = 32'd30
; 
32'd37692: dataIn1 = 32'd31
; 
32'd37693: dataIn1 = 32'd32
; 
32'd37694: dataIn1 = 32'd33
; 
32'd37695: dataIn1 = 32'd34
; 
32'd37696: dataIn1 = 32'd35
; 
32'd37697: dataIn1 = 32'd37
; 
32'd37698: dataIn1 = 32'd39
; 
32'd37699: dataIn1 = 32'd40
; 
32'd37700: dataIn1 = 32'd41
; 
32'd37701: dataIn1 = 32'd42
; 
32'd37702: dataIn1 = 32'd43
; 
32'd37703: dataIn1 = 32'd44
; 
32'd37704: dataIn1 = 32'd45
; 
32'd37705: dataIn1 = 32'd47
; 
32'd37706: dataIn1 = 32'd48
; 
32'd37707: dataIn1 = 32'd49
; 
32'd37708: dataIn1 = 32'd51
; 
32'd37709: dataIn1 = 32'd53
; 
32'd37710: dataIn1 = 32'd54
; 
32'd37711: dataIn1 = 32'd55
; 
32'd37712: dataIn1 = 32'd56
; 
32'd37713: dataIn1 = 32'd57
; 
32'd37714: dataIn1 = 32'd58
; 
32'd37715: dataIn1 = 32'd59
; 
32'd37716: dataIn1 = 32'd60
; 
32'd37717: dataIn1 = 32'd61
; 
32'd37718: dataIn1 = 32'd62
; 
32'd37719: dataIn1 = 32'd63
; 
32'd37720: dataIn1 = 32'd0
; 
32'd37721: dataIn1 = 32'd1
; 
32'd37722: dataIn1 = 32'd2
; 
32'd37723: dataIn1 = 32'd3
; 
32'd37724: dataIn1 = 32'd4
; 
32'd37725: dataIn1 = 32'd5
; 
32'd37726: dataIn1 = 32'd6
; 
32'd37727: dataIn1 = 32'd7
; 
32'd37728: dataIn1 = 32'd9
; 
32'd37729: dataIn1 = 32'd11
; 
32'd37730: dataIn1 = 32'd14
; 
32'd37731: dataIn1 = 32'd15
; 
32'd37732: dataIn1 = 32'd16
; 
32'd37733: dataIn1 = 32'd18
; 
32'd37734: dataIn1 = 32'd19
; 
32'd37735: dataIn1 = 32'd20
; 
32'd37736: dataIn1 = 32'd21
; 
32'd37737: dataIn1 = 32'd22
; 
32'd37738: dataIn1 = 32'd23
; 
32'd37739: dataIn1 = 32'd24
; 
32'd37740: dataIn1 = 32'd25
; 
32'd37741: dataIn1 = 32'd26
; 
32'd37742: dataIn1 = 32'd27
; 
32'd37743: dataIn1 = 32'd29
; 
32'd37744: dataIn1 = 32'd30
; 
32'd37745: dataIn1 = 32'd31
; 
32'd37746: dataIn1 = 32'd32
; 
32'd37747: dataIn1 = 32'd33
; 
32'd37748: dataIn1 = 32'd34
; 
32'd37749: dataIn1 = 32'd35
; 
32'd37750: dataIn1 = 32'd36
; 
32'd37751: dataIn1 = 32'd38
; 
32'd37752: dataIn1 = 32'd39
; 
32'd37753: dataIn1 = 32'd40
; 
32'd37754: dataIn1 = 32'd41
; 
32'd37755: dataIn1 = 32'd43
; 
32'd37756: dataIn1 = 32'd44
; 
32'd37757: dataIn1 = 32'd45
; 
32'd37758: dataIn1 = 32'd47
; 
32'd37759: dataIn1 = 32'd48
; 
32'd37760: dataIn1 = 32'd49
; 
32'd37761: dataIn1 = 32'd51
; 
32'd37762: dataIn1 = 32'd52
; 
32'd37763: dataIn1 = 32'd53
; 
32'd37764: dataIn1 = 32'd56
; 
32'd37765: dataIn1 = 32'd57
; 
32'd37766: dataIn1 = 32'd58
; 
32'd37767: dataIn1 = 32'd59
; 
32'd37768: dataIn1 = 32'd60
; 
32'd37769: dataIn1 = 32'd61
; 
32'd37770: dataIn1 = 32'd62
; 
32'd37771: dataIn1 = 32'd2
; 
32'd37772: dataIn1 = 32'd3
; 
32'd37773: dataIn1 = 32'd4
; 
32'd37774: dataIn1 = 32'd6
; 
32'd37775: dataIn1 = 32'd9
; 
32'd37776: dataIn1 = 32'd10
; 
32'd37777: dataIn1 = 32'd11
; 
32'd37778: dataIn1 = 32'd12
; 
32'd37779: dataIn1 = 32'd13
; 
32'd37780: dataIn1 = 32'd14
; 
32'd37781: dataIn1 = 32'd15
; 
32'd37782: dataIn1 = 32'd17
; 
32'd37783: dataIn1 = 32'd18
; 
32'd37784: dataIn1 = 32'd19
; 
32'd37785: dataIn1 = 32'd20
; 
32'd37786: dataIn1 = 32'd21
; 
32'd37787: dataIn1 = 32'd22
; 
32'd37788: dataIn1 = 32'd23
; 
32'd37789: dataIn1 = 32'd24
; 
32'd37790: dataIn1 = 32'd25
; 
32'd37791: dataIn1 = 32'd26
; 
32'd37792: dataIn1 = 32'd27
; 
32'd37793: dataIn1 = 32'd29
; 
32'd37794: dataIn1 = 32'd31
; 
32'd37795: dataIn1 = 32'd33
; 
32'd37796: dataIn1 = 32'd34
; 
32'd37797: dataIn1 = 32'd35
; 
32'd37798: dataIn1 = 32'd36
; 
32'd37799: dataIn1 = 32'd37
; 
32'd37800: dataIn1 = 32'd39
; 
32'd37801: dataIn1 = 32'd40
; 
32'd37802: dataIn1 = 32'd41
; 
32'd37803: dataIn1 = 32'd42
; 
32'd37804: dataIn1 = 32'd43
; 
32'd37805: dataIn1 = 32'd44
; 
32'd37806: dataIn1 = 32'd45
; 
32'd37807: dataIn1 = 32'd46
; 
32'd37808: dataIn1 = 32'd47
; 
32'd37809: dataIn1 = 32'd50
; 
32'd37810: dataIn1 = 32'd53
; 
32'd37811: dataIn1 = 32'd54
; 
32'd37812: dataIn1 = 32'd56
; 
32'd37813: dataIn1 = 32'd57
; 
32'd37814: dataIn1 = 32'd58
; 
32'd37815: dataIn1 = 32'd59
; 
32'd37816: dataIn1 = 32'd60
; 
32'd37817: dataIn1 = 32'd62
; 
32'd37818: dataIn1 = 32'd0
; 
32'd37819: dataIn1 = 32'd1
; 
32'd37820: dataIn1 = 32'd2
; 
32'd37821: dataIn1 = 32'd3
; 
32'd37822: dataIn1 = 32'd4
; 
32'd37823: dataIn1 = 32'd5
; 
32'd37824: dataIn1 = 32'd6
; 
32'd37825: dataIn1 = 32'd7
; 
32'd37826: dataIn1 = 32'd9
; 
32'd37827: dataIn1 = 32'd10
; 
32'd37828: dataIn1 = 32'd11
; 
32'd37829: dataIn1 = 32'd12
; 
32'd37830: dataIn1 = 32'd14
; 
32'd37831: dataIn1 = 32'd15
; 
32'd37832: dataIn1 = 32'd16
; 
32'd37833: dataIn1 = 32'd18
; 
32'd37834: dataIn1 = 32'd20
; 
32'd37835: dataIn1 = 32'd21
; 
32'd37836: dataIn1 = 32'd24
; 
32'd37837: dataIn1 = 32'd27
; 
32'd37838: dataIn1 = 32'd29
; 
32'd37839: dataIn1 = 32'd30
; 
32'd37840: dataIn1 = 32'd31
; 
32'd37841: dataIn1 = 32'd32
; 
32'd37842: dataIn1 = 32'd35
; 
32'd37843: dataIn1 = 32'd36
; 
32'd37844: dataIn1 = 32'd39
; 
32'd37845: dataIn1 = 32'd40
; 
32'd37846: dataIn1 = 32'd41
; 
32'd37847: dataIn1 = 32'd43
; 
32'd37848: dataIn1 = 32'd44
; 
32'd37849: dataIn1 = 32'd45
; 
32'd37850: dataIn1 = 32'd46
; 
32'd37851: dataIn1 = 32'd47
; 
32'd37852: dataIn1 = 32'd48
; 
32'd37853: dataIn1 = 32'd49
; 
32'd37854: dataIn1 = 32'd51
; 
32'd37855: dataIn1 = 32'd53
; 
32'd37856: dataIn1 = 32'd54
; 
32'd37857: dataIn1 = 32'd55
; 
32'd37858: dataIn1 = 32'd56
; 
32'd37859: dataIn1 = 32'd57
; 
32'd37860: dataIn1 = 32'd59
; 
32'd37861: dataIn1 = 32'd60
; 
32'd37862: dataIn1 = 32'd61
; 
32'd37863: dataIn1 = 32'd62
; 
32'd37864: dataIn1 = 32'd63
; 
32'd37865: dataIn1 = 32'd0
; 
32'd37866: dataIn1 = 32'd1
; 
32'd37867: dataIn1 = 32'd2
; 
32'd37868: dataIn1 = 32'd3
; 
32'd37869: dataIn1 = 32'd4
; 
32'd37870: dataIn1 = 32'd5
; 
32'd37871: dataIn1 = 32'd6
; 
32'd37872: dataIn1 = 32'd7
; 
32'd37873: dataIn1 = 32'd8
; 
32'd37874: dataIn1 = 32'd10
; 
32'd37875: dataIn1 = 32'd11
; 
32'd37876: dataIn1 = 32'd12
; 
32'd37877: dataIn1 = 32'd13
; 
32'd37878: dataIn1 = 32'd14
; 
32'd37879: dataIn1 = 32'd16
; 
32'd37880: dataIn1 = 32'd17
; 
32'd37881: dataIn1 = 32'd18
; 
32'd37882: dataIn1 = 32'd19
; 
32'd37883: dataIn1 = 32'd20
; 
32'd37884: dataIn1 = 32'd21
; 
32'd37885: dataIn1 = 32'd22
; 
32'd37886: dataIn1 = 32'd23
; 
32'd37887: dataIn1 = 32'd24
; 
32'd37888: dataIn1 = 32'd26
; 
32'd37889: dataIn1 = 32'd27
; 
32'd37890: dataIn1 = 32'd28
; 
32'd37891: dataIn1 = 32'd31
; 
32'd37892: dataIn1 = 32'd33
; 
32'd37893: dataIn1 = 32'd35
; 
32'd37894: dataIn1 = 32'd36
; 
32'd37895: dataIn1 = 32'd37
; 
32'd37896: dataIn1 = 32'd38
; 
32'd37897: dataIn1 = 32'd39
; 
32'd37898: dataIn1 = 32'd40
; 
32'd37899: dataIn1 = 32'd42
; 
32'd37900: dataIn1 = 32'd44
; 
32'd37901: dataIn1 = 32'd45
; 
32'd37902: dataIn1 = 32'd46
; 
32'd37903: dataIn1 = 32'd47
; 
32'd37904: dataIn1 = 32'd48
; 
32'd37905: dataIn1 = 32'd49
; 
32'd37906: dataIn1 = 32'd50
; 
32'd37907: dataIn1 = 32'd51
; 
32'd37908: dataIn1 = 32'd52
; 
32'd37909: dataIn1 = 32'd53
; 
32'd37910: dataIn1 = 32'd54
; 
32'd37911: dataIn1 = 32'd55
; 
32'd37912: dataIn1 = 32'd57
; 
32'd37913: dataIn1 = 32'd58
; 
32'd37914: dataIn1 = 32'd59
; 
32'd37915: dataIn1 = 32'd60
; 
32'd37916: dataIn1 = 32'd61
; 
32'd37917: dataIn1 = 32'd62
; 
32'd37918: dataIn1 = 32'd63
; 
32'd37919: dataIn1 = 32'd0
; 
32'd37920: dataIn1 = 32'd1
; 
32'd37921: dataIn1 = 32'd2
; 
32'd37922: dataIn1 = 32'd3
; 
32'd37923: dataIn1 = 32'd4
; 
32'd37924: dataIn1 = 32'd5
; 
32'd37925: dataIn1 = 32'd6
; 
32'd37926: dataIn1 = 32'd7
; 
32'd37927: dataIn1 = 32'd8
; 
32'd37928: dataIn1 = 32'd9
; 
32'd37929: dataIn1 = 32'd10
; 
32'd37930: dataIn1 = 32'd11
; 
32'd37931: dataIn1 = 32'd12
; 
32'd37932: dataIn1 = 32'd13
; 
32'd37933: dataIn1 = 32'd14
; 
32'd37934: dataIn1 = 32'd15
; 
32'd37935: dataIn1 = 32'd16
; 
32'd37936: dataIn1 = 32'd17
; 
32'd37937: dataIn1 = 32'd18
; 
32'd37938: dataIn1 = 32'd19
; 
32'd37939: dataIn1 = 32'd21
; 
32'd37940: dataIn1 = 32'd22
; 
32'd37941: dataIn1 = 32'd23
; 
32'd37942: dataIn1 = 32'd24
; 
32'd37943: dataIn1 = 32'd25
; 
32'd37944: dataIn1 = 32'd27
; 
32'd37945: dataIn1 = 32'd28
; 
32'd37946: dataIn1 = 32'd29
; 
32'd37947: dataIn1 = 32'd30
; 
32'd37948: dataIn1 = 32'd31
; 
32'd37949: dataIn1 = 32'd33
; 
32'd37950: dataIn1 = 32'd34
; 
32'd37951: dataIn1 = 32'd35
; 
32'd37952: dataIn1 = 32'd38
; 
32'd37953: dataIn1 = 32'd39
; 
32'd37954: dataIn1 = 32'd40
; 
32'd37955: dataIn1 = 32'd41
; 
32'd37956: dataIn1 = 32'd42
; 
32'd37957: dataIn1 = 32'd43
; 
32'd37958: dataIn1 = 32'd45
; 
32'd37959: dataIn1 = 32'd46
; 
32'd37960: dataIn1 = 32'd47
; 
32'd37961: dataIn1 = 32'd48
; 
32'd37962: dataIn1 = 32'd50
; 
32'd37963: dataIn1 = 32'd51
; 
32'd37964: dataIn1 = 32'd52
; 
32'd37965: dataIn1 = 32'd54
; 
32'd37966: dataIn1 = 32'd55
; 
32'd37967: dataIn1 = 32'd56
; 
32'd37968: dataIn1 = 32'd57
; 
32'd37969: dataIn1 = 32'd59
; 
32'd37970: dataIn1 = 32'd60
; 
32'd37971: dataIn1 = 32'd61
; 
32'd37972: dataIn1 = 32'd63
; 
32'd37973: dataIn1 = 32'd0
; 
32'd37974: dataIn1 = 32'd2
; 
32'd37975: dataIn1 = 32'd4
; 
32'd37976: dataIn1 = 32'd5
; 
32'd37977: dataIn1 = 32'd6
; 
32'd37978: dataIn1 = 32'd7
; 
32'd37979: dataIn1 = 32'd10
; 
32'd37980: dataIn1 = 32'd11
; 
32'd37981: dataIn1 = 32'd14
; 
32'd37982: dataIn1 = 32'd16
; 
32'd37983: dataIn1 = 32'd17
; 
32'd37984: dataIn1 = 32'd18
; 
32'd37985: dataIn1 = 32'd21
; 
32'd37986: dataIn1 = 32'd22
; 
32'd37987: dataIn1 = 32'd23
; 
32'd37988: dataIn1 = 32'd25
; 
32'd37989: dataIn1 = 32'd26
; 
32'd37990: dataIn1 = 32'd27
; 
32'd37991: dataIn1 = 32'd29
; 
32'd37992: dataIn1 = 32'd30
; 
32'd37993: dataIn1 = 32'd31
; 
32'd37994: dataIn1 = 32'd32
; 
32'd37995: dataIn1 = 32'd33
; 
32'd37996: dataIn1 = 32'd34
; 
32'd37997: dataIn1 = 32'd35
; 
32'd37998: dataIn1 = 32'd36
; 
32'd37999: dataIn1 = 32'd37
; 
32'd38000: dataIn1 = 32'd38
; 
32'd38001: dataIn1 = 32'd39
; 
32'd38002: dataIn1 = 32'd40
; 
32'd38003: dataIn1 = 32'd42
; 
32'd38004: dataIn1 = 32'd43
; 
32'd38005: dataIn1 = 32'd44
; 
32'd38006: dataIn1 = 32'd45
; 
32'd38007: dataIn1 = 32'd46
; 
32'd38008: dataIn1 = 32'd47
; 
32'd38009: dataIn1 = 32'd48
; 
32'd38010: dataIn1 = 32'd50
; 
32'd38011: dataIn1 = 32'd53
; 
32'd38012: dataIn1 = 32'd54
; 
32'd38013: dataIn1 = 32'd55
; 
32'd38014: dataIn1 = 32'd56
; 
32'd38015: dataIn1 = 32'd57
; 
32'd38016: dataIn1 = 32'd59
; 
32'd38017: dataIn1 = 32'd61
; 
32'd38018: dataIn1 = 32'd62
; 
32'd38019: dataIn1 = 32'd63
; 
32'd38020: dataIn1 = 32'd0
; 
32'd38021: dataIn1 = 32'd1
; 
32'd38022: dataIn1 = 32'd2
; 
32'd38023: dataIn1 = 32'd3
; 
32'd38024: dataIn1 = 32'd5
; 
32'd38025: dataIn1 = 32'd6
; 
32'd38026: dataIn1 = 32'd7
; 
32'd38027: dataIn1 = 32'd8
; 
32'd38028: dataIn1 = 32'd9
; 
32'd38029: dataIn1 = 32'd10
; 
32'd38030: dataIn1 = 32'd11
; 
32'd38031: dataIn1 = 32'd12
; 
32'd38032: dataIn1 = 32'd13
; 
32'd38033: dataIn1 = 32'd14
; 
32'd38034: dataIn1 = 32'd15
; 
32'd38035: dataIn1 = 32'd16
; 
32'd38036: dataIn1 = 32'd19
; 
32'd38037: dataIn1 = 32'd20
; 
32'd38038: dataIn1 = 32'd21
; 
32'd38039: dataIn1 = 32'd22
; 
32'd38040: dataIn1 = 32'd23
; 
32'd38041: dataIn1 = 32'd24
; 
32'd38042: dataIn1 = 32'd25
; 
32'd38043: dataIn1 = 32'd27
; 
32'd38044: dataIn1 = 32'd28
; 
32'd38045: dataIn1 = 32'd29
; 
32'd38046: dataIn1 = 32'd30
; 
32'd38047: dataIn1 = 32'd31
; 
32'd38048: dataIn1 = 32'd32
; 
32'd38049: dataIn1 = 32'd33
; 
32'd38050: dataIn1 = 32'd35
; 
32'd38051: dataIn1 = 32'd36
; 
32'd38052: dataIn1 = 32'd37
; 
32'd38053: dataIn1 = 32'd38
; 
32'd38054: dataIn1 = 32'd39
; 
32'd38055: dataIn1 = 32'd41
; 
32'd38056: dataIn1 = 32'd45
; 
32'd38057: dataIn1 = 32'd46
; 
32'd38058: dataIn1 = 32'd48
; 
32'd38059: dataIn1 = 32'd50
; 
32'd38060: dataIn1 = 32'd51
; 
32'd38061: dataIn1 = 32'd52
; 
32'd38062: dataIn1 = 32'd53
; 
32'd38063: dataIn1 = 32'd54
; 
32'd38064: dataIn1 = 32'd55
; 
32'd38065: dataIn1 = 32'd56
; 
32'd38066: dataIn1 = 32'd57
; 
32'd38067: dataIn1 = 32'd58
; 
32'd38068: dataIn1 = 32'd60
; 
32'd38069: dataIn1 = 32'd61
; 
32'd38070: dataIn1 = 32'd62
; 
32'd38071: dataIn1 = 32'd0
; 
32'd38072: dataIn1 = 32'd1
; 
32'd38073: dataIn1 = 32'd3
; 
32'd38074: dataIn1 = 32'd4
; 
32'd38075: dataIn1 = 32'd5
; 
32'd38076: dataIn1 = 32'd6
; 
32'd38077: dataIn1 = 32'd7
; 
32'd38078: dataIn1 = 32'd9
; 
32'd38079: dataIn1 = 32'd10
; 
32'd38080: dataIn1 = 32'd11
; 
32'd38081: dataIn1 = 32'd12
; 
32'd38082: dataIn1 = 32'd14
; 
32'd38083: dataIn1 = 32'd15
; 
32'd38084: dataIn1 = 32'd17
; 
32'd38085: dataIn1 = 32'd18
; 
32'd38086: dataIn1 = 32'd19
; 
32'd38087: dataIn1 = 32'd20
; 
32'd38088: dataIn1 = 32'd21
; 
32'd38089: dataIn1 = 32'd23
; 
32'd38090: dataIn1 = 32'd24
; 
32'd38091: dataIn1 = 32'd28
; 
32'd38092: dataIn1 = 32'd29
; 
32'd38093: dataIn1 = 32'd30
; 
32'd38094: dataIn1 = 32'd31
; 
32'd38095: dataIn1 = 32'd32
; 
32'd38096: dataIn1 = 32'd33
; 
32'd38097: dataIn1 = 32'd34
; 
32'd38098: dataIn1 = 32'd35
; 
32'd38099: dataIn1 = 32'd37
; 
32'd38100: dataIn1 = 32'd38
; 
32'd38101: dataIn1 = 32'd39
; 
32'd38102: dataIn1 = 32'd41
; 
32'd38103: dataIn1 = 32'd42
; 
32'd38104: dataIn1 = 32'd43
; 
32'd38105: dataIn1 = 32'd45
; 
32'd38106: dataIn1 = 32'd47
; 
32'd38107: dataIn1 = 32'd48
; 
32'd38108: dataIn1 = 32'd49
; 
32'd38109: dataIn1 = 32'd51
; 
32'd38110: dataIn1 = 32'd52
; 
32'd38111: dataIn1 = 32'd53
; 
32'd38112: dataIn1 = 32'd54
; 
32'd38113: dataIn1 = 32'd56
; 
32'd38114: dataIn1 = 32'd57
; 
32'd38115: dataIn1 = 32'd58
; 
32'd38116: dataIn1 = 32'd59
; 
32'd38117: dataIn1 = 32'd61
; 
32'd38118: dataIn1 = 32'd63
; 
32'd38119: dataIn1 = 32'd1
; 
32'd38120: dataIn1 = 32'd2
; 
32'd38121: dataIn1 = 32'd5
; 
32'd38122: dataIn1 = 32'd6
; 
32'd38123: dataIn1 = 32'd7
; 
32'd38124: dataIn1 = 32'd8
; 
32'd38125: dataIn1 = 32'd9
; 
32'd38126: dataIn1 = 32'd10
; 
32'd38127: dataIn1 = 32'd11
; 
32'd38128: dataIn1 = 32'd12
; 
32'd38129: dataIn1 = 32'd13
; 
32'd38130: dataIn1 = 32'd15
; 
32'd38131: dataIn1 = 32'd16
; 
32'd38132: dataIn1 = 32'd17
; 
32'd38133: dataIn1 = 32'd18
; 
32'd38134: dataIn1 = 32'd19
; 
32'd38135: dataIn1 = 32'd23
; 
32'd38136: dataIn1 = 32'd24
; 
32'd38137: dataIn1 = 32'd25
; 
32'd38138: dataIn1 = 32'd26
; 
32'd38139: dataIn1 = 32'd28
; 
32'd38140: dataIn1 = 32'd31
; 
32'd38141: dataIn1 = 32'd33
; 
32'd38142: dataIn1 = 32'd34
; 
32'd38143: dataIn1 = 32'd35
; 
32'd38144: dataIn1 = 32'd36
; 
32'd38145: dataIn1 = 32'd38
; 
32'd38146: dataIn1 = 32'd40
; 
32'd38147: dataIn1 = 32'd41
; 
32'd38148: dataIn1 = 32'd43
; 
32'd38149: dataIn1 = 32'd44
; 
32'd38150: dataIn1 = 32'd45
; 
32'd38151: dataIn1 = 32'd46
; 
32'd38152: dataIn1 = 32'd47
; 
32'd38153: dataIn1 = 32'd48
; 
32'd38154: dataIn1 = 32'd49
; 
32'd38155: dataIn1 = 32'd51
; 
32'd38156: dataIn1 = 32'd52
; 
32'd38157: dataIn1 = 32'd53
; 
32'd38158: dataIn1 = 32'd54
; 
32'd38159: dataIn1 = 32'd56
; 
32'd38160: dataIn1 = 32'd57
; 
32'd38161: dataIn1 = 32'd58
; 
32'd38162: dataIn1 = 32'd59
; 
32'd38163: dataIn1 = 32'd60
; 
32'd38164: dataIn1 = 32'd61
; 
32'd38165: dataIn1 = 32'd62
; 
32'd38166: dataIn1 = 32'd63
; 
32'd38167: dataIn1 = 32'd0
; 
32'd38168: dataIn1 = 32'd1
; 
32'd38169: dataIn1 = 32'd2
; 
32'd38170: dataIn1 = 32'd3
; 
32'd38171: dataIn1 = 32'd4
; 
32'd38172: dataIn1 = 32'd5
; 
32'd38173: dataIn1 = 32'd6
; 
32'd38174: dataIn1 = 32'd7
; 
32'd38175: dataIn1 = 32'd8
; 
32'd38176: dataIn1 = 32'd9
; 
32'd38177: dataIn1 = 32'd10
; 
32'd38178: dataIn1 = 32'd11
; 
32'd38179: dataIn1 = 32'd12
; 
32'd38180: dataIn1 = 32'd13
; 
32'd38181: dataIn1 = 32'd14
; 
32'd38182: dataIn1 = 32'd15
; 
32'd38183: dataIn1 = 32'd16
; 
32'd38184: dataIn1 = 32'd18
; 
32'd38185: dataIn1 = 32'd19
; 
32'd38186: dataIn1 = 32'd20
; 
32'd38187: dataIn1 = 32'd21
; 
32'd38188: dataIn1 = 32'd22
; 
32'd38189: dataIn1 = 32'd24
; 
32'd38190: dataIn1 = 32'd26
; 
32'd38191: dataIn1 = 32'd27
; 
32'd38192: dataIn1 = 32'd28
; 
32'd38193: dataIn1 = 32'd29
; 
32'd38194: dataIn1 = 32'd30
; 
32'd38195: dataIn1 = 32'd32
; 
32'd38196: dataIn1 = 32'd34
; 
32'd38197: dataIn1 = 32'd35
; 
32'd38198: dataIn1 = 32'd36
; 
32'd38199: dataIn1 = 32'd37
; 
32'd38200: dataIn1 = 32'd38
; 
32'd38201: dataIn1 = 32'd39
; 
32'd38202: dataIn1 = 32'd41
; 
32'd38203: dataIn1 = 32'd42
; 
32'd38204: dataIn1 = 32'd43
; 
32'd38205: dataIn1 = 32'd44
; 
32'd38206: dataIn1 = 32'd45
; 
32'd38207: dataIn1 = 32'd47
; 
32'd38208: dataIn1 = 32'd48
; 
32'd38209: dataIn1 = 32'd49
; 
32'd38210: dataIn1 = 32'd50
; 
32'd38211: dataIn1 = 32'd51
; 
32'd38212: dataIn1 = 32'd52
; 
32'd38213: dataIn1 = 32'd53
; 
32'd38214: dataIn1 = 32'd55
; 
32'd38215: dataIn1 = 32'd56
; 
32'd38216: dataIn1 = 32'd58
; 
32'd38217: dataIn1 = 32'd59
; 
32'd38218: dataIn1 = 32'd61
; 
32'd38219: dataIn1 = 32'd62
; 
32'd38220: dataIn1 = 32'd63
; 
32'd38221: dataIn1 = 32'd0
; 
32'd38222: dataIn1 = 32'd2
; 
32'd38223: dataIn1 = 32'd3
; 
32'd38224: dataIn1 = 32'd4
; 
32'd38225: dataIn1 = 32'd5
; 
32'd38226: dataIn1 = 32'd6
; 
32'd38227: dataIn1 = 32'd7
; 
32'd38228: dataIn1 = 32'd8
; 
32'd38229: dataIn1 = 32'd9
; 
32'd38230: dataIn1 = 32'd10
; 
32'd38231: dataIn1 = 32'd11
; 
32'd38232: dataIn1 = 32'd12
; 
32'd38233: dataIn1 = 32'd13
; 
32'd38234: dataIn1 = 32'd14
; 
32'd38235: dataIn1 = 32'd15
; 
32'd38236: dataIn1 = 32'd16
; 
32'd38237: dataIn1 = 32'd18
; 
32'd38238: dataIn1 = 32'd19
; 
32'd38239: dataIn1 = 32'd20
; 
32'd38240: dataIn1 = 32'd21
; 
32'd38241: dataIn1 = 32'd22
; 
32'd38242: dataIn1 = 32'd23
; 
32'd38243: dataIn1 = 32'd24
; 
32'd38244: dataIn1 = 32'd25
; 
32'd38245: dataIn1 = 32'd27
; 
32'd38246: dataIn1 = 32'd28
; 
32'd38247: dataIn1 = 32'd29
; 
32'd38248: dataIn1 = 32'd30
; 
32'd38249: dataIn1 = 32'd32
; 
32'd38250: dataIn1 = 32'd33
; 
32'd38251: dataIn1 = 32'd35
; 
32'd38252: dataIn1 = 32'd36
; 
32'd38253: dataIn1 = 32'd37
; 
32'd38254: dataIn1 = 32'd38
; 
32'd38255: dataIn1 = 32'd39
; 
32'd38256: dataIn1 = 32'd40
; 
32'd38257: dataIn1 = 32'd41
; 
32'd38258: dataIn1 = 32'd42
; 
32'd38259: dataIn1 = 32'd43
; 
32'd38260: dataIn1 = 32'd44
; 
32'd38261: dataIn1 = 32'd45
; 
32'd38262: dataIn1 = 32'd47
; 
32'd38263: dataIn1 = 32'd50
; 
32'd38264: dataIn1 = 32'd53
; 
32'd38265: dataIn1 = 32'd54
; 
32'd38266: dataIn1 = 32'd55
; 
32'd38267: dataIn1 = 32'd57
; 
32'd38268: dataIn1 = 32'd59
; 
32'd38269: dataIn1 = 32'd60
; 
32'd38270: dataIn1 = 32'd61
; 
32'd38271: dataIn1 = 32'd62
; 
32'd38272: dataIn1 = 32'd63
; 
32'd38273: dataIn1 = 32'd0
; 
32'd38274: dataIn1 = 32'd1
; 
32'd38275: dataIn1 = 32'd2
; 
32'd38276: dataIn1 = 32'd3
; 
32'd38277: dataIn1 = 32'd5
; 
32'd38278: dataIn1 = 32'd8
; 
32'd38279: dataIn1 = 32'd9
; 
32'd38280: dataIn1 = 32'd10
; 
32'd38281: dataIn1 = 32'd12
; 
32'd38282: dataIn1 = 32'd13
; 
32'd38283: dataIn1 = 32'd14
; 
32'd38284: dataIn1 = 32'd15
; 
32'd38285: dataIn1 = 32'd16
; 
32'd38286: dataIn1 = 32'd17
; 
32'd38287: dataIn1 = 32'd21
; 
32'd38288: dataIn1 = 32'd22
; 
32'd38289: dataIn1 = 32'd23
; 
32'd38290: dataIn1 = 32'd25
; 
32'd38291: dataIn1 = 32'd27
; 
32'd38292: dataIn1 = 32'd28
; 
32'd38293: dataIn1 = 32'd29
; 
32'd38294: dataIn1 = 32'd30
; 
32'd38295: dataIn1 = 32'd32
; 
32'd38296: dataIn1 = 32'd33
; 
32'd38297: dataIn1 = 32'd34
; 
32'd38298: dataIn1 = 32'd35
; 
32'd38299: dataIn1 = 32'd37
; 
32'd38300: dataIn1 = 32'd38
; 
32'd38301: dataIn1 = 32'd40
; 
32'd38302: dataIn1 = 32'd41
; 
32'd38303: dataIn1 = 32'd42
; 
32'd38304: dataIn1 = 32'd43
; 
32'd38305: dataIn1 = 32'd44
; 
32'd38306: dataIn1 = 32'd45
; 
32'd38307: dataIn1 = 32'd46
; 
32'd38308: dataIn1 = 32'd48
; 
32'd38309: dataIn1 = 32'd49
; 
32'd38310: dataIn1 = 32'd50
; 
32'd38311: dataIn1 = 32'd51
; 
32'd38312: dataIn1 = 32'd52
; 
32'd38313: dataIn1 = 32'd53
; 
32'd38314: dataIn1 = 32'd54
; 
32'd38315: dataIn1 = 32'd55
; 
32'd38316: dataIn1 = 32'd57
; 
32'd38317: dataIn1 = 32'd58
; 
32'd38318: dataIn1 = 32'd59
; 
32'd38319: dataIn1 = 32'd60
; 
32'd38320: dataIn1 = 32'd61
; 
32'd38321: dataIn1 = 32'd63
; 
32'd38322: dataIn1 = 32'd0
; 
32'd38323: dataIn1 = 32'd1
; 
32'd38324: dataIn1 = 32'd3
; 
32'd38325: dataIn1 = 32'd4
; 
32'd38326: dataIn1 = 32'd5
; 
32'd38327: dataIn1 = 32'd6
; 
32'd38328: dataIn1 = 32'd7
; 
32'd38329: dataIn1 = 32'd8
; 
32'd38330: dataIn1 = 32'd10
; 
32'd38331: dataIn1 = 32'd12
; 
32'd38332: dataIn1 = 32'd14
; 
32'd38333: dataIn1 = 32'd16
; 
32'd38334: dataIn1 = 32'd18
; 
32'd38335: dataIn1 = 32'd21
; 
32'd38336: dataIn1 = 32'd24
; 
32'd38337: dataIn1 = 32'd25
; 
32'd38338: dataIn1 = 32'd26
; 
32'd38339: dataIn1 = 32'd27
; 
32'd38340: dataIn1 = 32'd28
; 
32'd38341: dataIn1 = 32'd30
; 
32'd38342: dataIn1 = 32'd31
; 
32'd38343: dataIn1 = 32'd33
; 
32'd38344: dataIn1 = 32'd34
; 
32'd38345: dataIn1 = 32'd35
; 
32'd38346: dataIn1 = 32'd36
; 
32'd38347: dataIn1 = 32'd37
; 
32'd38348: dataIn1 = 32'd38
; 
32'd38349: dataIn1 = 32'd39
; 
32'd38350: dataIn1 = 32'd40
; 
32'd38351: dataIn1 = 32'd42
; 
32'd38352: dataIn1 = 32'd43
; 
32'd38353: dataIn1 = 32'd44
; 
32'd38354: dataIn1 = 32'd46
; 
32'd38355: dataIn1 = 32'd47
; 
32'd38356: dataIn1 = 32'd48
; 
32'd38357: dataIn1 = 32'd49
; 
32'd38358: dataIn1 = 32'd50
; 
32'd38359: dataIn1 = 32'd52
; 
32'd38360: dataIn1 = 32'd53
; 
32'd38361: dataIn1 = 32'd54
; 
32'd38362: dataIn1 = 32'd57
; 
32'd38363: dataIn1 = 32'd58
; 
32'd38364: dataIn1 = 32'd59
; 
32'd38365: dataIn1 = 32'd60
; 
32'd38366: dataIn1 = 32'd61
; 
32'd38367: dataIn1 = 32'd62
; 
32'd38368: dataIn1 = 32'd63
; 
32'd38369: dataIn1 = 32'd1
; 
32'd38370: dataIn1 = 32'd3
; 
32'd38371: dataIn1 = 32'd4
; 
32'd38372: dataIn1 = 32'd5
; 
32'd38373: dataIn1 = 32'd6
; 
32'd38374: dataIn1 = 32'd7
; 
32'd38375: dataIn1 = 32'd8
; 
32'd38376: dataIn1 = 32'd9
; 
32'd38377: dataIn1 = 32'd10
; 
32'd38378: dataIn1 = 32'd12
; 
32'd38379: dataIn1 = 32'd13
; 
32'd38380: dataIn1 = 32'd14
; 
32'd38381: dataIn1 = 32'd16
; 
32'd38382: dataIn1 = 32'd17
; 
32'd38383: dataIn1 = 32'd18
; 
32'd38384: dataIn1 = 32'd19
; 
32'd38385: dataIn1 = 32'd20
; 
32'd38386: dataIn1 = 32'd21
; 
32'd38387: dataIn1 = 32'd22
; 
32'd38388: dataIn1 = 32'd24
; 
32'd38389: dataIn1 = 32'd25
; 
32'd38390: dataIn1 = 32'd29
; 
32'd38391: dataIn1 = 32'd30
; 
32'd38392: dataIn1 = 32'd31
; 
32'd38393: dataIn1 = 32'd32
; 
32'd38394: dataIn1 = 32'd33
; 
32'd38395: dataIn1 = 32'd34
; 
32'd38396: dataIn1 = 32'd38
; 
32'd38397: dataIn1 = 32'd40
; 
32'd38398: dataIn1 = 32'd42
; 
32'd38399: dataIn1 = 32'd44
; 
32'd38400: dataIn1 = 32'd45
; 
32'd38401: dataIn1 = 32'd46
; 
32'd38402: dataIn1 = 32'd47
; 
32'd38403: dataIn1 = 32'd48
; 
32'd38404: dataIn1 = 32'd49
; 
32'd38405: dataIn1 = 32'd50
; 
32'd38406: dataIn1 = 32'd51
; 
32'd38407: dataIn1 = 32'd53
; 
32'd38408: dataIn1 = 32'd54
; 
32'd38409: dataIn1 = 32'd55
; 
32'd38410: dataIn1 = 32'd57
; 
32'd38411: dataIn1 = 32'd58
; 
32'd38412: dataIn1 = 32'd60
; 
32'd38413: dataIn1 = 32'd61
; 
32'd38414: dataIn1 = 32'd62
; 
32'd38415: dataIn1 = 32'd0
; 
32'd38416: dataIn1 = 32'd1
; 
32'd38417: dataIn1 = 32'd2
; 
32'd38418: dataIn1 = 32'd3
; 
32'd38419: dataIn1 = 32'd4
; 
32'd38420: dataIn1 = 32'd6
; 
32'd38421: dataIn1 = 32'd7
; 
32'd38422: dataIn1 = 32'd8
; 
32'd38423: dataIn1 = 32'd9
; 
32'd38424: dataIn1 = 32'd10
; 
32'd38425: dataIn1 = 32'd12
; 
32'd38426: dataIn1 = 32'd13
; 
32'd38427: dataIn1 = 32'd15
; 
32'd38428: dataIn1 = 32'd16
; 
32'd38429: dataIn1 = 32'd17
; 
32'd38430: dataIn1 = 32'd19
; 
32'd38431: dataIn1 = 32'd20
; 
32'd38432: dataIn1 = 32'd21
; 
32'd38433: dataIn1 = 32'd22
; 
32'd38434: dataIn1 = 32'd24
; 
32'd38435: dataIn1 = 32'd25
; 
32'd38436: dataIn1 = 32'd27
; 
32'd38437: dataIn1 = 32'd28
; 
32'd38438: dataIn1 = 32'd29
; 
32'd38439: dataIn1 = 32'd30
; 
32'd38440: dataIn1 = 32'd32
; 
32'd38441: dataIn1 = 32'd33
; 
32'd38442: dataIn1 = 32'd34
; 
32'd38443: dataIn1 = 32'd35
; 
32'd38444: dataIn1 = 32'd36
; 
32'd38445: dataIn1 = 32'd37
; 
32'd38446: dataIn1 = 32'd38
; 
32'd38447: dataIn1 = 32'd39
; 
32'd38448: dataIn1 = 32'd41
; 
32'd38449: dataIn1 = 32'd42
; 
32'd38450: dataIn1 = 32'd43
; 
32'd38451: dataIn1 = 32'd45
; 
32'd38452: dataIn1 = 32'd47
; 
32'd38453: dataIn1 = 32'd48
; 
32'd38454: dataIn1 = 32'd49
; 
32'd38455: dataIn1 = 32'd51
; 
32'd38456: dataIn1 = 32'd52
; 
32'd38457: dataIn1 = 32'd53
; 
32'd38458: dataIn1 = 32'd54
; 
32'd38459: dataIn1 = 32'd55
; 
32'd38460: dataIn1 = 32'd56
; 
32'd38461: dataIn1 = 32'd58
; 
32'd38462: dataIn1 = 32'd59
; 
32'd38463: dataIn1 = 32'd61
; 
32'd38464: dataIn1 = 32'd62
; 
32'd38465: dataIn1 = 32'd63
; 
32'd38466: dataIn1 = 32'd0
; 
32'd38467: dataIn1 = 32'd2
; 
32'd38468: dataIn1 = 32'd3
; 
32'd38469: dataIn1 = 32'd4
; 
32'd38470: dataIn1 = 32'd5
; 
32'd38471: dataIn1 = 32'd6
; 
32'd38472: dataIn1 = 32'd7
; 
32'd38473: dataIn1 = 32'd8
; 
32'd38474: dataIn1 = 32'd9
; 
32'd38475: dataIn1 = 32'd10
; 
32'd38476: dataIn1 = 32'd11
; 
32'd38477: dataIn1 = 32'd13
; 
32'd38478: dataIn1 = 32'd14
; 
32'd38479: dataIn1 = 32'd15
; 
32'd38480: dataIn1 = 32'd16
; 
32'd38481: dataIn1 = 32'd17
; 
32'd38482: dataIn1 = 32'd18
; 
32'd38483: dataIn1 = 32'd19
; 
32'd38484: dataIn1 = 32'd21
; 
32'd38485: dataIn1 = 32'd24
; 
32'd38486: dataIn1 = 32'd25
; 
32'd38487: dataIn1 = 32'd26
; 
32'd38488: dataIn1 = 32'd27
; 
32'd38489: dataIn1 = 32'd28
; 
32'd38490: dataIn1 = 32'd30
; 
32'd38491: dataIn1 = 32'd31
; 
32'd38492: dataIn1 = 32'd33
; 
32'd38493: dataIn1 = 32'd35
; 
32'd38494: dataIn1 = 32'd37
; 
32'd38495: dataIn1 = 32'd38
; 
32'd38496: dataIn1 = 32'd39
; 
32'd38497: dataIn1 = 32'd41
; 
32'd38498: dataIn1 = 32'd42
; 
32'd38499: dataIn1 = 32'd43
; 
32'd38500: dataIn1 = 32'd44
; 
32'd38501: dataIn1 = 32'd45
; 
32'd38502: dataIn1 = 32'd46
; 
32'd38503: dataIn1 = 32'd47
; 
32'd38504: dataIn1 = 32'd48
; 
32'd38505: dataIn1 = 32'd49
; 
32'd38506: dataIn1 = 32'd50
; 
32'd38507: dataIn1 = 32'd51
; 
32'd38508: dataIn1 = 32'd52
; 
32'd38509: dataIn1 = 32'd53
; 
32'd38510: dataIn1 = 32'd54
; 
32'd38511: dataIn1 = 32'd55
; 
32'd38512: dataIn1 = 32'd56
; 
32'd38513: dataIn1 = 32'd57
; 
32'd38514: dataIn1 = 32'd59
; 
32'd38515: dataIn1 = 32'd60
; 
32'd38516: dataIn1 = 32'd61
; 
32'd38517: dataIn1 = 32'd62
; 
32'd38518: dataIn1 = 32'd63
; 
32'd38519: dataIn1 = 32'd0
; 
32'd38520: dataIn1 = 32'd2
; 
32'd38521: dataIn1 = 32'd7
; 
32'd38522: dataIn1 = 32'd8
; 
32'd38523: dataIn1 = 32'd9
; 
32'd38524: dataIn1 = 32'd10
; 
32'd38525: dataIn1 = 32'd11
; 
32'd38526: dataIn1 = 32'd12
; 
32'd38527: dataIn1 = 32'd13
; 
32'd38528: dataIn1 = 32'd16
; 
32'd38529: dataIn1 = 32'd17
; 
32'd38530: dataIn1 = 32'd18
; 
32'd38531: dataIn1 = 32'd19
; 
32'd38532: dataIn1 = 32'd20
; 
32'd38533: dataIn1 = 32'd21
; 
32'd38534: dataIn1 = 32'd22
; 
32'd38535: dataIn1 = 32'd23
; 
32'd38536: dataIn1 = 32'd24
; 
32'd38537: dataIn1 = 32'd25
; 
32'd38538: dataIn1 = 32'd26
; 
32'd38539: dataIn1 = 32'd27
; 
32'd38540: dataIn1 = 32'd28
; 
32'd38541: dataIn1 = 32'd29
; 
32'd38542: dataIn1 = 32'd30
; 
32'd38543: dataIn1 = 32'd31
; 
32'd38544: dataIn1 = 32'd32
; 
32'd38545: dataIn1 = 32'd33
; 
32'd38546: dataIn1 = 32'd35
; 
32'd38547: dataIn1 = 32'd36
; 
32'd38548: dataIn1 = 32'd38
; 
32'd38549: dataIn1 = 32'd40
; 
32'd38550: dataIn1 = 32'd41
; 
32'd38551: dataIn1 = 32'd42
; 
32'd38552: dataIn1 = 32'd43
; 
32'd38553: dataIn1 = 32'd44
; 
32'd38554: dataIn1 = 32'd46
; 
32'd38555: dataIn1 = 32'd47
; 
32'd38556: dataIn1 = 32'd50
; 
32'd38557: dataIn1 = 32'd51
; 
32'd38558: dataIn1 = 32'd53
; 
32'd38559: dataIn1 = 32'd54
; 
32'd38560: dataIn1 = 32'd55
; 
32'd38561: dataIn1 = 32'd56
; 
32'd38562: dataIn1 = 32'd57
; 
32'd38563: dataIn1 = 32'd59
; 
32'd38564: dataIn1 = 32'd60
; 
32'd38565: dataIn1 = 32'd61
; 
32'd38566: dataIn1 = 32'd63
; 
32'd38567: dataIn1 = 32'd0
; 
32'd38568: dataIn1 = 32'd4
; 
32'd38569: dataIn1 = 32'd5
; 
32'd38570: dataIn1 = 32'd6
; 
32'd38571: dataIn1 = 32'd7
; 
32'd38572: dataIn1 = 32'd8
; 
32'd38573: dataIn1 = 32'd9
; 
32'd38574: dataIn1 = 32'd11
; 
32'd38575: dataIn1 = 32'd13
; 
32'd38576: dataIn1 = 32'd14
; 
32'd38577: dataIn1 = 32'd15
; 
32'd38578: dataIn1 = 32'd16
; 
32'd38579: dataIn1 = 32'd17
; 
32'd38580: dataIn1 = 32'd18
; 
32'd38581: dataIn1 = 32'd19
; 
32'd38582: dataIn1 = 32'd20
; 
32'd38583: dataIn1 = 32'd21
; 
32'd38584: dataIn1 = 32'd22
; 
32'd38585: dataIn1 = 32'd23
; 
32'd38586: dataIn1 = 32'd24
; 
32'd38587: dataIn1 = 32'd25
; 
32'd38588: dataIn1 = 32'd26
; 
32'd38589: dataIn1 = 32'd30
; 
32'd38590: dataIn1 = 32'd31
; 
32'd38591: dataIn1 = 32'd32
; 
32'd38592: dataIn1 = 32'd33
; 
32'd38593: dataIn1 = 32'd34
; 
32'd38594: dataIn1 = 32'd36
; 
32'd38595: dataIn1 = 32'd37
; 
32'd38596: dataIn1 = 32'd38
; 
32'd38597: dataIn1 = 32'd40
; 
32'd38598: dataIn1 = 32'd41
; 
32'd38599: dataIn1 = 32'd42
; 
32'd38600: dataIn1 = 32'd43
; 
32'd38601: dataIn1 = 32'd45
; 
32'd38602: dataIn1 = 32'd46
; 
32'd38603: dataIn1 = 32'd47
; 
32'd38604: dataIn1 = 32'd48
; 
32'd38605: dataIn1 = 32'd51
; 
32'd38606: dataIn1 = 32'd53
; 
32'd38607: dataIn1 = 32'd54
; 
32'd38608: dataIn1 = 32'd55
; 
32'd38609: dataIn1 = 32'd56
; 
32'd38610: dataIn1 = 32'd57
; 
32'd38611: dataIn1 = 32'd59
; 
32'd38612: dataIn1 = 32'd60
; 
32'd38613: dataIn1 = 32'd61
; 
32'd38614: dataIn1 = 32'd62
; 
32'd38615: dataIn1 = 32'd0
; 
32'd38616: dataIn1 = 32'd1
; 
32'd38617: dataIn1 = 32'd3
; 
32'd38618: dataIn1 = 32'd4
; 
32'd38619: dataIn1 = 32'd6
; 
32'd38620: dataIn1 = 32'd7
; 
32'd38621: dataIn1 = 32'd8
; 
32'd38622: dataIn1 = 32'd9
; 
32'd38623: dataIn1 = 32'd10
; 
32'd38624: dataIn1 = 32'd11
; 
32'd38625: dataIn1 = 32'd12
; 
32'd38626: dataIn1 = 32'd13
; 
32'd38627: dataIn1 = 32'd15
; 
32'd38628: dataIn1 = 32'd16
; 
32'd38629: dataIn1 = 32'd17
; 
32'd38630: dataIn1 = 32'd19
; 
32'd38631: dataIn1 = 32'd20
; 
32'd38632: dataIn1 = 32'd23
; 
32'd38633: dataIn1 = 32'd27
; 
32'd38634: dataIn1 = 32'd30
; 
32'd38635: dataIn1 = 32'd31
; 
32'd38636: dataIn1 = 32'd32
; 
32'd38637: dataIn1 = 32'd33
; 
32'd38638: dataIn1 = 32'd35
; 
32'd38639: dataIn1 = 32'd36
; 
32'd38640: dataIn1 = 32'd37
; 
32'd38641: dataIn1 = 32'd38
; 
32'd38642: dataIn1 = 32'd41
; 
32'd38643: dataIn1 = 32'd42
; 
32'd38644: dataIn1 = 32'd43
; 
32'd38645: dataIn1 = 32'd44
; 
32'd38646: dataIn1 = 32'd45
; 
32'd38647: dataIn1 = 32'd46
; 
32'd38648: dataIn1 = 32'd47
; 
32'd38649: dataIn1 = 32'd48
; 
32'd38650: dataIn1 = 32'd50
; 
32'd38651: dataIn1 = 32'd51
; 
32'd38652: dataIn1 = 32'd52
; 
32'd38653: dataIn1 = 32'd53
; 
32'd38654: dataIn1 = 32'd54
; 
32'd38655: dataIn1 = 32'd55
; 
32'd38656: dataIn1 = 32'd56
; 
32'd38657: dataIn1 = 32'd58
; 
32'd38658: dataIn1 = 32'd59
; 
32'd38659: dataIn1 = 32'd61
; 
32'd38660: dataIn1 = 32'd63
; 
32'd38661: dataIn1 = 32'd0
; 
32'd38662: dataIn1 = 32'd1
; 
32'd38663: dataIn1 = 32'd2
; 
32'd38664: dataIn1 = 32'd3
; 
32'd38665: dataIn1 = 32'd4
; 
32'd38666: dataIn1 = 32'd5
; 
32'd38667: dataIn1 = 32'd7
; 
32'd38668: dataIn1 = 32'd8
; 
32'd38669: dataIn1 = 32'd10
; 
32'd38670: dataIn1 = 32'd11
; 
32'd38671: dataIn1 = 32'd12
; 
32'd38672: dataIn1 = 32'd14
; 
32'd38673: dataIn1 = 32'd15
; 
32'd38674: dataIn1 = 32'd16
; 
32'd38675: dataIn1 = 32'd18
; 
32'd38676: dataIn1 = 32'd19
; 
32'd38677: dataIn1 = 32'd20
; 
32'd38678: dataIn1 = 32'd21
; 
32'd38679: dataIn1 = 32'd22
; 
32'd38680: dataIn1 = 32'd23
; 
32'd38681: dataIn1 = 32'd24
; 
32'd38682: dataIn1 = 32'd25
; 
32'd38683: dataIn1 = 32'd26
; 
32'd38684: dataIn1 = 32'd29
; 
32'd38685: dataIn1 = 32'd30
; 
32'd38686: dataIn1 = 32'd32
; 
32'd38687: dataIn1 = 32'd33
; 
32'd38688: dataIn1 = 32'd34
; 
32'd38689: dataIn1 = 32'd35
; 
32'd38690: dataIn1 = 32'd36
; 
32'd38691: dataIn1 = 32'd37
; 
32'd38692: dataIn1 = 32'd39
; 
32'd38693: dataIn1 = 32'd40
; 
32'd38694: dataIn1 = 32'd41
; 
32'd38695: dataIn1 = 32'd43
; 
32'd38696: dataIn1 = 32'd44
; 
32'd38697: dataIn1 = 32'd46
; 
32'd38698: dataIn1 = 32'd47
; 
32'd38699: dataIn1 = 32'd48
; 
32'd38700: dataIn1 = 32'd49
; 
32'd38701: dataIn1 = 32'd52
; 
32'd38702: dataIn1 = 32'd54
; 
32'd38703: dataIn1 = 32'd55
; 
32'd38704: dataIn1 = 32'd56
; 
32'd38705: dataIn1 = 32'd59
; 
32'd38706: dataIn1 = 32'd60
; 
32'd38707: dataIn1 = 32'd62
; 
32'd38708: dataIn1 = 32'd63
; 
32'd38709: dataIn1 = 32'd0
; 
32'd38710: dataIn1 = 32'd1
; 
32'd38711: dataIn1 = 32'd2
; 
32'd38712: dataIn1 = 32'd3
; 
32'd38713: dataIn1 = 32'd4
; 
32'd38714: dataIn1 = 32'd5
; 
32'd38715: dataIn1 = 32'd6
; 
32'd38716: dataIn1 = 32'd7
; 
32'd38717: dataIn1 = 32'd9
; 
32'd38718: dataIn1 = 32'd10
; 
32'd38719: dataIn1 = 32'd12
; 
32'd38720: dataIn1 = 32'd13
; 
32'd38721: dataIn1 = 32'd14
; 
32'd38722: dataIn1 = 32'd15
; 
32'd38723: dataIn1 = 32'd16
; 
32'd38724: dataIn1 = 32'd17
; 
32'd38725: dataIn1 = 32'd18
; 
32'd38726: dataIn1 = 32'd21
; 
32'd38727: dataIn1 = 32'd22
; 
32'd38728: dataIn1 = 32'd23
; 
32'd38729: dataIn1 = 32'd24
; 
32'd38730: dataIn1 = 32'd25
; 
32'd38731: dataIn1 = 32'd26
; 
32'd38732: dataIn1 = 32'd27
; 
32'd38733: dataIn1 = 32'd28
; 
32'd38734: dataIn1 = 32'd29
; 
32'd38735: dataIn1 = 32'd30
; 
32'd38736: dataIn1 = 32'd31
; 
32'd38737: dataIn1 = 32'd32
; 
32'd38738: dataIn1 = 32'd33
; 
32'd38739: dataIn1 = 32'd35
; 
32'd38740: dataIn1 = 32'd36
; 
32'd38741: dataIn1 = 32'd37
; 
32'd38742: dataIn1 = 32'd40
; 
32'd38743: dataIn1 = 32'd41
; 
32'd38744: dataIn1 = 32'd44
; 
32'd38745: dataIn1 = 32'd45
; 
32'd38746: dataIn1 = 32'd47
; 
32'd38747: dataIn1 = 32'd48
; 
32'd38748: dataIn1 = 32'd49
; 
32'd38749: dataIn1 = 32'd51
; 
32'd38750: dataIn1 = 32'd52
; 
32'd38751: dataIn1 = 32'd53
; 
32'd38752: dataIn1 = 32'd54
; 
32'd38753: dataIn1 = 32'd55
; 
32'd38754: dataIn1 = 32'd57
; 
32'd38755: dataIn1 = 32'd58
; 
32'd38756: dataIn1 = 32'd60
; 
32'd38757: dataIn1 = 32'd61
; 
32'd38758: dataIn1 = 32'd62
; 
32'd38759: dataIn1 = 32'd63
; 
32'd38760: dataIn1 = 32'd0
; 
32'd38761: dataIn1 = 32'd2
; 
32'd38762: dataIn1 = 32'd3
; 
32'd38763: dataIn1 = 32'd4
; 
32'd38764: dataIn1 = 32'd5
; 
32'd38765: dataIn1 = 32'd6
; 
32'd38766: dataIn1 = 32'd8
; 
32'd38767: dataIn1 = 32'd9
; 
32'd38768: dataIn1 = 32'd12
; 
32'd38769: dataIn1 = 32'd13
; 
32'd38770: dataIn1 = 32'd14
; 
32'd38771: dataIn1 = 32'd15
; 
32'd38772: dataIn1 = 32'd17
; 
32'd38773: dataIn1 = 32'd18
; 
32'd38774: dataIn1 = 32'd19
; 
32'd38775: dataIn1 = 32'd20
; 
32'd38776: dataIn1 = 32'd21
; 
32'd38777: dataIn1 = 32'd22
; 
32'd38778: dataIn1 = 32'd23
; 
32'd38779: dataIn1 = 32'd24
; 
32'd38780: dataIn1 = 32'd25
; 
32'd38781: dataIn1 = 32'd26
; 
32'd38782: dataIn1 = 32'd27
; 
32'd38783: dataIn1 = 32'd28
; 
32'd38784: dataIn1 = 32'd29
; 
32'd38785: dataIn1 = 32'd30
; 
32'd38786: dataIn1 = 32'd31
; 
32'd38787: dataIn1 = 32'd33
; 
32'd38788: dataIn1 = 32'd35
; 
32'd38789: dataIn1 = 32'd36
; 
32'd38790: dataIn1 = 32'd37
; 
32'd38791: dataIn1 = 32'd38
; 
32'd38792: dataIn1 = 32'd39
; 
32'd38793: dataIn1 = 32'd41
; 
32'd38794: dataIn1 = 32'd42
; 
32'd38795: dataIn1 = 32'd44
; 
32'd38796: dataIn1 = 32'd45
; 
32'd38797: dataIn1 = 32'd46
; 
32'd38798: dataIn1 = 32'd47
; 
32'd38799: dataIn1 = 32'd48
; 
32'd38800: dataIn1 = 32'd50
; 
32'd38801: dataIn1 = 32'd51
; 
32'd38802: dataIn1 = 32'd53
; 
32'd38803: dataIn1 = 32'd54
; 
32'd38804: dataIn1 = 32'd55
; 
32'd38805: dataIn1 = 32'd56
; 
32'd38806: dataIn1 = 32'd57
; 
32'd38807: dataIn1 = 32'd58
; 
32'd38808: dataIn1 = 32'd59
; 
32'd38809: dataIn1 = 32'd60
; 
32'd38810: dataIn1 = 32'd62
; 
32'd38811: dataIn1 = 32'd0
; 
32'd38812: dataIn1 = 32'd1
; 
32'd38813: dataIn1 = 32'd2
; 
32'd38814: dataIn1 = 32'd3
; 
32'd38815: dataIn1 = 32'd4
; 
32'd38816: dataIn1 = 32'd5
; 
32'd38817: dataIn1 = 32'd6
; 
32'd38818: dataIn1 = 32'd7
; 
32'd38819: dataIn1 = 32'd10
; 
32'd38820: dataIn1 = 32'd11
; 
32'd38821: dataIn1 = 32'd12
; 
32'd38822: dataIn1 = 32'd13
; 
32'd38823: dataIn1 = 32'd14
; 
32'd38824: dataIn1 = 32'd15
; 
32'd38825: dataIn1 = 32'd16
; 
32'd38826: dataIn1 = 32'd18
; 
32'd38827: dataIn1 = 32'd19
; 
32'd38828: dataIn1 = 32'd20
; 
32'd38829: dataIn1 = 32'd21
; 
32'd38830: dataIn1 = 32'd22
; 
32'd38831: dataIn1 = 32'd23
; 
32'd38832: dataIn1 = 32'd25
; 
32'd38833: dataIn1 = 32'd27
; 
32'd38834: dataIn1 = 32'd28
; 
32'd38835: dataIn1 = 32'd29
; 
32'd38836: dataIn1 = 32'd30
; 
32'd38837: dataIn1 = 32'd31
; 
32'd38838: dataIn1 = 32'd32
; 
32'd38839: dataIn1 = 32'd34
; 
32'd38840: dataIn1 = 32'd35
; 
32'd38841: dataIn1 = 32'd36
; 
32'd38842: dataIn1 = 32'd38
; 
32'd38843: dataIn1 = 32'd39
; 
32'd38844: dataIn1 = 32'd40
; 
32'd38845: dataIn1 = 32'd41
; 
32'd38846: dataIn1 = 32'd42
; 
32'd38847: dataIn1 = 32'd43
; 
32'd38848: dataIn1 = 32'd45
; 
32'd38849: dataIn1 = 32'd46
; 
32'd38850: dataIn1 = 32'd47
; 
32'd38851: dataIn1 = 32'd49
; 
32'd38852: dataIn1 = 32'd50
; 
32'd38853: dataIn1 = 32'd51
; 
32'd38854: dataIn1 = 32'd53
; 
32'd38855: dataIn1 = 32'd54
; 
32'd38856: dataIn1 = 32'd55
; 
32'd38857: dataIn1 = 32'd57
; 
32'd38858: dataIn1 = 32'd58
; 
32'd38859: dataIn1 = 32'd59
; 
32'd38860: dataIn1 = 32'd60
; 
32'd38861: dataIn1 = 32'd61
; 
32'd38862: dataIn1 = 32'd63
; 
32'd38863: dataIn1 = 32'd1
; 
32'd38864: dataIn1 = 32'd2
; 
32'd38865: dataIn1 = 32'd3
; 
32'd38866: dataIn1 = 32'd4
; 
32'd38867: dataIn1 = 32'd5
; 
32'd38868: dataIn1 = 32'd6
; 
32'd38869: dataIn1 = 32'd7
; 
32'd38870: dataIn1 = 32'd10
; 
32'd38871: dataIn1 = 32'd11
; 
32'd38872: dataIn1 = 32'd12
; 
32'd38873: dataIn1 = 32'd13
; 
32'd38874: dataIn1 = 32'd14
; 
32'd38875: dataIn1 = 32'd16
; 
32'd38876: dataIn1 = 32'd17
; 
32'd38877: dataIn1 = 32'd18
; 
32'd38878: dataIn1 = 32'd20
; 
32'd38879: dataIn1 = 32'd22
; 
32'd38880: dataIn1 = 32'd23
; 
32'd38881: dataIn1 = 32'd24
; 
32'd38882: dataIn1 = 32'd25
; 
32'd38883: dataIn1 = 32'd26
; 
32'd38884: dataIn1 = 32'd27
; 
32'd38885: dataIn1 = 32'd28
; 
32'd38886: dataIn1 = 32'd29
; 
32'd38887: dataIn1 = 32'd30
; 
32'd38888: dataIn1 = 32'd31
; 
32'd38889: dataIn1 = 32'd32
; 
32'd38890: dataIn1 = 32'd33
; 
32'd38891: dataIn1 = 32'd34
; 
32'd38892: dataIn1 = 32'd35
; 
32'd38893: dataIn1 = 32'd36
; 
32'd38894: dataIn1 = 32'd37
; 
32'd38895: dataIn1 = 32'd38
; 
32'd38896: dataIn1 = 32'd39
; 
32'd38897: dataIn1 = 32'd40
; 
32'd38898: dataIn1 = 32'd43
; 
32'd38899: dataIn1 = 32'd44
; 
32'd38900: dataIn1 = 32'd46
; 
32'd38901: dataIn1 = 32'd47
; 
32'd38902: dataIn1 = 32'd48
; 
32'd38903: dataIn1 = 32'd50
; 
32'd38904: dataIn1 = 32'd53
; 
32'd38905: dataIn1 = 32'd55
; 
32'd38906: dataIn1 = 32'd56
; 
32'd38907: dataIn1 = 32'd57
; 
32'd38908: dataIn1 = 32'd58
; 
32'd38909: dataIn1 = 32'd59
; 
32'd38910: dataIn1 = 32'd60
; 
32'd38911: dataIn1 = 32'd61
; 
32'd38912: dataIn1 = 32'd62
; 
32'd38913: dataIn1 = 32'd63
; 
32'd38914: dataIn1 = 32'd0
; 
32'd38915: dataIn1 = 32'd1
; 
32'd38916: dataIn1 = 32'd2
; 
32'd38917: dataIn1 = 32'd5
; 
32'd38918: dataIn1 = 32'd6
; 
32'd38919: dataIn1 = 32'd7
; 
32'd38920: dataIn1 = 32'd8
; 
32'd38921: dataIn1 = 32'd9
; 
32'd38922: dataIn1 = 32'd10
; 
32'd38923: dataIn1 = 32'd11
; 
32'd38924: dataIn1 = 32'd12
; 
32'd38925: dataIn1 = 32'd13
; 
32'd38926: dataIn1 = 32'd14
; 
32'd38927: dataIn1 = 32'd15
; 
32'd38928: dataIn1 = 32'd16
; 
32'd38929: dataIn1 = 32'd17
; 
32'd38930: dataIn1 = 32'd18
; 
32'd38931: dataIn1 = 32'd19
; 
32'd38932: dataIn1 = 32'd21
; 
32'd38933: dataIn1 = 32'd22
; 
32'd38934: dataIn1 = 32'd23
; 
32'd38935: dataIn1 = 32'd24
; 
32'd38936: dataIn1 = 32'd26
; 
32'd38937: dataIn1 = 32'd27
; 
32'd38938: dataIn1 = 32'd29
; 
32'd38939: dataIn1 = 32'd31
; 
32'd38940: dataIn1 = 32'd33
; 
32'd38941: dataIn1 = 32'd35
; 
32'd38942: dataIn1 = 32'd36
; 
32'd38943: dataIn1 = 32'd37
; 
32'd38944: dataIn1 = 32'd38
; 
32'd38945: dataIn1 = 32'd40
; 
32'd38946: dataIn1 = 32'd42
; 
32'd38947: dataIn1 = 32'd44
; 
32'd38948: dataIn1 = 32'd45
; 
32'd38949: dataIn1 = 32'd47
; 
32'd38950: dataIn1 = 32'd48
; 
32'd38951: dataIn1 = 32'd49
; 
32'd38952: dataIn1 = 32'd50
; 
32'd38953: dataIn1 = 32'd52
; 
32'd38954: dataIn1 = 32'd54
; 
32'd38955: dataIn1 = 32'd55
; 
32'd38956: dataIn1 = 32'd56
; 
32'd38957: dataIn1 = 32'd57
; 
32'd38958: dataIn1 = 32'd58
; 
32'd38959: dataIn1 = 32'd59
; 
32'd38960: dataIn1 = 32'd60
; 
32'd38961: dataIn1 = 32'd61
; 
32'd38962: dataIn1 = 32'd62
; 
32'd38963: dataIn1 = 32'd63
; 
32'd38964: dataIn1 = 32'd1
; 
32'd38965: dataIn1 = 32'd2
; 
32'd38966: dataIn1 = 32'd3
; 
32'd38967: dataIn1 = 32'd5
; 
32'd38968: dataIn1 = 32'd6
; 
32'd38969: dataIn1 = 32'd7
; 
32'd38970: dataIn1 = 32'd9
; 
32'd38971: dataIn1 = 32'd11
; 
32'd38972: dataIn1 = 32'd12
; 
32'd38973: dataIn1 = 32'd13
; 
32'd38974: dataIn1 = 32'd14
; 
32'd38975: dataIn1 = 32'd15
; 
32'd38976: dataIn1 = 32'd16
; 
32'd38977: dataIn1 = 32'd17
; 
32'd38978: dataIn1 = 32'd18
; 
32'd38979: dataIn1 = 32'd19
; 
32'd38980: dataIn1 = 32'd20
; 
32'd38981: dataIn1 = 32'd21
; 
32'd38982: dataIn1 = 32'd22
; 
32'd38983: dataIn1 = 32'd25
; 
32'd38984: dataIn1 = 32'd27
; 
32'd38985: dataIn1 = 32'd29
; 
32'd38986: dataIn1 = 32'd30
; 
32'd38987: dataIn1 = 32'd32
; 
32'd38988: dataIn1 = 32'd34
; 
32'd38989: dataIn1 = 32'd35
; 
32'd38990: dataIn1 = 32'd36
; 
32'd38991: dataIn1 = 32'd37
; 
32'd38992: dataIn1 = 32'd38
; 
32'd38993: dataIn1 = 32'd39
; 
32'd38994: dataIn1 = 32'd40
; 
32'd38995: dataIn1 = 32'd41
; 
32'd38996: dataIn1 = 32'd42
; 
32'd38997: dataIn1 = 32'd43
; 
32'd38998: dataIn1 = 32'd44
; 
32'd38999: dataIn1 = 32'd45
; 
32'd39000: dataIn1 = 32'd47
; 
32'd39001: dataIn1 = 32'd48
; 
32'd39002: dataIn1 = 32'd50
; 
32'd39003: dataIn1 = 32'd51
; 
32'd39004: dataIn1 = 32'd53
; 
32'd39005: dataIn1 = 32'd55
; 
32'd39006: dataIn1 = 32'd57
; 
32'd39007: dataIn1 = 32'd58
; 
32'd39008: dataIn1 = 32'd59
; 
32'd39009: dataIn1 = 32'd61
; 
32'd39010: dataIn1 = 32'd62
; 
32'd39011: dataIn1 = 32'd63
; 
32'd39012: dataIn1 = 32'd1
; 
32'd39013: dataIn1 = 32'd2
; 
32'd39014: dataIn1 = 32'd4
; 
32'd39015: dataIn1 = 32'd5
; 
32'd39016: dataIn1 = 32'd7
; 
32'd39017: dataIn1 = 32'd8
; 
32'd39018: dataIn1 = 32'd9
; 
32'd39019: dataIn1 = 32'd10
; 
32'd39020: dataIn1 = 32'd11
; 
32'd39021: dataIn1 = 32'd12
; 
32'd39022: dataIn1 = 32'd13
; 
32'd39023: dataIn1 = 32'd16
; 
32'd39024: dataIn1 = 32'd18
; 
32'd39025: dataIn1 = 32'd19
; 
32'd39026: dataIn1 = 32'd20
; 
32'd39027: dataIn1 = 32'd22
; 
32'd39028: dataIn1 = 32'd23
; 
32'd39029: dataIn1 = 32'd24
; 
32'd39030: dataIn1 = 32'd25
; 
32'd39031: dataIn1 = 32'd26
; 
32'd39032: dataIn1 = 32'd27
; 
32'd39033: dataIn1 = 32'd28
; 
32'd39034: dataIn1 = 32'd29
; 
32'd39035: dataIn1 = 32'd30
; 
32'd39036: dataIn1 = 32'd31
; 
32'd39037: dataIn1 = 32'd32
; 
32'd39038: dataIn1 = 32'd34
; 
32'd39039: dataIn1 = 32'd35
; 
32'd39040: dataIn1 = 32'd36
; 
32'd39041: dataIn1 = 32'd38
; 
32'd39042: dataIn1 = 32'd42
; 
32'd39043: dataIn1 = 32'd43
; 
32'd39044: dataIn1 = 32'd44
; 
32'd39045: dataIn1 = 32'd45
; 
32'd39046: dataIn1 = 32'd46
; 
32'd39047: dataIn1 = 32'd47
; 
32'd39048: dataIn1 = 32'd48
; 
32'd39049: dataIn1 = 32'd49
; 
32'd39050: dataIn1 = 32'd50
; 
32'd39051: dataIn1 = 32'd51
; 
32'd39052: dataIn1 = 32'd52
; 
32'd39053: dataIn1 = 32'd53
; 
32'd39054: dataIn1 = 32'd54
; 
32'd39055: dataIn1 = 32'd56
; 
32'd39056: dataIn1 = 32'd57
; 
32'd39057: dataIn1 = 32'd58
; 
32'd39058: dataIn1 = 32'd59
; 
32'd39059: dataIn1 = 32'd60
; 
32'd39060: dataIn1 = 32'd61
; 
32'd39061: dataIn1 = 32'd62
; 
32'd39062: dataIn1 = 32'd63
; 
32'd39063: dataIn1 = 32'd0
; 
32'd39064: dataIn1 = 32'd1
; 
32'd39065: dataIn1 = 32'd2
; 
32'd39066: dataIn1 = 32'd3
; 
32'd39067: dataIn1 = 32'd4
; 
32'd39068: dataIn1 = 32'd5
; 
32'd39069: dataIn1 = 32'd6
; 
32'd39070: dataIn1 = 32'd7
; 
32'd39071: dataIn1 = 32'd8
; 
32'd39072: dataIn1 = 32'd9
; 
32'd39073: dataIn1 = 32'd11
; 
32'd39074: dataIn1 = 32'd12
; 
32'd39075: dataIn1 = 32'd13
; 
32'd39076: dataIn1 = 32'd14
; 
32'd39077: dataIn1 = 32'd15
; 
32'd39078: dataIn1 = 32'd16
; 
32'd39079: dataIn1 = 32'd17
; 
32'd39080: dataIn1 = 32'd18
; 
32'd39081: dataIn1 = 32'd20
; 
32'd39082: dataIn1 = 32'd22
; 
32'd39083: dataIn1 = 32'd23
; 
32'd39084: dataIn1 = 32'd25
; 
32'd39085: dataIn1 = 32'd26
; 
32'd39086: dataIn1 = 32'd28
; 
32'd39087: dataIn1 = 32'd29
; 
32'd39088: dataIn1 = 32'd30
; 
32'd39089: dataIn1 = 32'd31
; 
32'd39090: dataIn1 = 32'd32
; 
32'd39091: dataIn1 = 32'd33
; 
32'd39092: dataIn1 = 32'd34
; 
32'd39093: dataIn1 = 32'd36
; 
32'd39094: dataIn1 = 32'd38
; 
32'd39095: dataIn1 = 32'd39
; 
32'd39096: dataIn1 = 32'd41
; 
32'd39097: dataIn1 = 32'd42
; 
32'd39098: dataIn1 = 32'd43
; 
32'd39099: dataIn1 = 32'd44
; 
32'd39100: dataIn1 = 32'd45
; 
32'd39101: dataIn1 = 32'd46
; 
32'd39102: dataIn1 = 32'd48
; 
32'd39103: dataIn1 = 32'd49
; 
32'd39104: dataIn1 = 32'd50
; 
32'd39105: dataIn1 = 32'd51
; 
32'd39106: dataIn1 = 32'd52
; 
32'd39107: dataIn1 = 32'd53
; 
32'd39108: dataIn1 = 32'd54
; 
32'd39109: dataIn1 = 32'd55
; 
32'd39110: dataIn1 = 32'd56
; 
32'd39111: dataIn1 = 32'd58
; 
32'd39112: dataIn1 = 32'd59
; 
32'd39113: dataIn1 = 32'd63
; 
32'd39114: dataIn1 = 32'd0
; 
32'd39115: dataIn1 = 32'd1
; 
32'd39116: dataIn1 = 32'd3
; 
32'd39117: dataIn1 = 32'd4
; 
32'd39118: dataIn1 = 32'd5
; 
32'd39119: dataIn1 = 32'd6
; 
32'd39120: dataIn1 = 32'd7
; 
32'd39121: dataIn1 = 32'd9
; 
32'd39122: dataIn1 = 32'd10
; 
32'd39123: dataIn1 = 32'd11
; 
32'd39124: dataIn1 = 32'd12
; 
32'd39125: dataIn1 = 32'd13
; 
32'd39126: dataIn1 = 32'd14
; 
32'd39127: dataIn1 = 32'd15
; 
32'd39128: dataIn1 = 32'd16
; 
32'd39129: dataIn1 = 32'd17
; 
32'd39130: dataIn1 = 32'd18
; 
32'd39131: dataIn1 = 32'd19
; 
32'd39132: dataIn1 = 32'd20
; 
32'd39133: dataIn1 = 32'd21
; 
32'd39134: dataIn1 = 32'd22
; 
32'd39135: dataIn1 = 32'd23
; 
32'd39136: dataIn1 = 32'd24
; 
32'd39137: dataIn1 = 32'd26
; 
32'd39138: dataIn1 = 32'd28
; 
32'd39139: dataIn1 = 32'd29
; 
32'd39140: dataIn1 = 32'd31
; 
32'd39141: dataIn1 = 32'd32
; 
32'd39142: dataIn1 = 32'd35
; 
32'd39143: dataIn1 = 32'd36
; 
32'd39144: dataIn1 = 32'd37
; 
32'd39145: dataIn1 = 32'd38
; 
32'd39146: dataIn1 = 32'd40
; 
32'd39147: dataIn1 = 32'd43
; 
32'd39148: dataIn1 = 32'd45
; 
32'd39149: dataIn1 = 32'd46
; 
32'd39150: dataIn1 = 32'd48
; 
32'd39151: dataIn1 = 32'd49
; 
32'd39152: dataIn1 = 32'd50
; 
32'd39153: dataIn1 = 32'd51
; 
32'd39154: dataIn1 = 32'd53
; 
32'd39155: dataIn1 = 32'd54
; 
32'd39156: dataIn1 = 32'd58
; 
32'd39157: dataIn1 = 32'd59
; 
32'd39158: dataIn1 = 32'd60
; 
32'd39159: dataIn1 = 32'd61
; 
32'd39160: dataIn1 = 32'd63
; 
32'd39161: dataIn1 = 32'd0
; 
32'd39162: dataIn1 = 32'd2
; 
32'd39163: dataIn1 = 32'd3
; 
32'd39164: dataIn1 = 32'd5
; 
32'd39165: dataIn1 = 32'd6
; 
32'd39166: dataIn1 = 32'd7
; 
32'd39167: dataIn1 = 32'd8
; 
32'd39168: dataIn1 = 32'd9
; 
32'd39169: dataIn1 = 32'd10
; 
32'd39170: dataIn1 = 32'd12
; 
32'd39171: dataIn1 = 32'd13
; 
32'd39172: dataIn1 = 32'd14
; 
32'd39173: dataIn1 = 32'd15
; 
32'd39174: dataIn1 = 32'd16
; 
32'd39175: dataIn1 = 32'd17
; 
32'd39176: dataIn1 = 32'd18
; 
32'd39177: dataIn1 = 32'd19
; 
32'd39178: dataIn1 = 32'd20
; 
32'd39179: dataIn1 = 32'd21
; 
32'd39180: dataIn1 = 32'd22
; 
32'd39181: dataIn1 = 32'd23
; 
32'd39182: dataIn1 = 32'd24
; 
32'd39183: dataIn1 = 32'd27
; 
32'd39184: dataIn1 = 32'd28
; 
32'd39185: dataIn1 = 32'd32
; 
32'd39186: dataIn1 = 32'd33
; 
32'd39187: dataIn1 = 32'd34
; 
32'd39188: dataIn1 = 32'd35
; 
32'd39189: dataIn1 = 32'd36
; 
32'd39190: dataIn1 = 32'd38
; 
32'd39191: dataIn1 = 32'd39
; 
32'd39192: dataIn1 = 32'd40
; 
32'd39193: dataIn1 = 32'd41
; 
32'd39194: dataIn1 = 32'd42
; 
32'd39195: dataIn1 = 32'd43
; 
32'd39196: dataIn1 = 32'd44
; 
32'd39197: dataIn1 = 32'd46
; 
32'd39198: dataIn1 = 32'd48
; 
32'd39199: dataIn1 = 32'd49
; 
32'd39200: dataIn1 = 32'd50
; 
32'd39201: dataIn1 = 32'd52
; 
32'd39202: dataIn1 = 32'd53
; 
32'd39203: dataIn1 = 32'd54
; 
32'd39204: dataIn1 = 32'd55
; 
32'd39205: dataIn1 = 32'd56
; 
32'd39206: dataIn1 = 32'd58
; 
32'd39207: dataIn1 = 32'd59
; 
32'd39208: dataIn1 = 32'd61
; 
32'd39209: dataIn1 = 32'd62
; 
32'd39210: dataIn1 = 32'd63
; 
32'd39211: dataIn1 = 32'd0
; 
32'd39212: dataIn1 = 32'd2
; 
32'd39213: dataIn1 = 32'd4
; 
32'd39214: dataIn1 = 32'd5
; 
32'd39215: dataIn1 = 32'd6
; 
32'd39216: dataIn1 = 32'd7
; 
32'd39217: dataIn1 = 32'd8
; 
32'd39218: dataIn1 = 32'd9
; 
32'd39219: dataIn1 = 32'd11
; 
32'd39220: dataIn1 = 32'd12
; 
32'd39221: dataIn1 = 32'd13
; 
32'd39222: dataIn1 = 32'd14
; 
32'd39223: dataIn1 = 32'd16
; 
32'd39224: dataIn1 = 32'd17
; 
32'd39225: dataIn1 = 32'd21
; 
32'd39226: dataIn1 = 32'd22
; 
32'd39227: dataIn1 = 32'd24
; 
32'd39228: dataIn1 = 32'd26
; 
32'd39229: dataIn1 = 32'd27
; 
32'd39230: dataIn1 = 32'd29
; 
32'd39231: dataIn1 = 32'd30
; 
32'd39232: dataIn1 = 32'd31
; 
32'd39233: dataIn1 = 32'd33
; 
32'd39234: dataIn1 = 32'd35
; 
32'd39235: dataIn1 = 32'd37
; 
32'd39236: dataIn1 = 32'd38
; 
32'd39237: dataIn1 = 32'd39
; 
32'd39238: dataIn1 = 32'd40
; 
32'd39239: dataIn1 = 32'd43
; 
32'd39240: dataIn1 = 32'd45
; 
32'd39241: dataIn1 = 32'd46
; 
32'd39242: dataIn1 = 32'd50
; 
32'd39243: dataIn1 = 32'd51
; 
32'd39244: dataIn1 = 32'd54
; 
32'd39245: dataIn1 = 32'd55
; 
32'd39246: dataIn1 = 32'd56
; 
32'd39247: dataIn1 = 32'd57
; 
32'd39248: dataIn1 = 32'd58
; 
32'd39249: dataIn1 = 32'd59
; 
32'd39250: dataIn1 = 32'd60
; 
32'd39251: dataIn1 = 32'd61
; 
32'd39252: dataIn1 = 32'd62
; 
32'd39253: dataIn1 = 32'd1
; 
32'd39254: dataIn1 = 32'd2
; 
32'd39255: dataIn1 = 32'd4
; 
32'd39256: dataIn1 = 32'd5
; 
32'd39257: dataIn1 = 32'd6
; 
32'd39258: dataIn1 = 32'd8
; 
32'd39259: dataIn1 = 32'd9
; 
32'd39260: dataIn1 = 32'd10
; 
32'd39261: dataIn1 = 32'd11
; 
32'd39262: dataIn1 = 32'd12
; 
32'd39263: dataIn1 = 32'd13
; 
32'd39264: dataIn1 = 32'd14
; 
32'd39265: dataIn1 = 32'd15
; 
32'd39266: dataIn1 = 32'd16
; 
32'd39267: dataIn1 = 32'd18
; 
32'd39268: dataIn1 = 32'd19
; 
32'd39269: dataIn1 = 32'd21
; 
32'd39270: dataIn1 = 32'd22
; 
32'd39271: dataIn1 = 32'd23
; 
32'd39272: dataIn1 = 32'd25
; 
32'd39273: dataIn1 = 32'd26
; 
32'd39274: dataIn1 = 32'd27
; 
32'd39275: dataIn1 = 32'd30
; 
32'd39276: dataIn1 = 32'd31
; 
32'd39277: dataIn1 = 32'd33
; 
32'd39278: dataIn1 = 32'd34
; 
32'd39279: dataIn1 = 32'd35
; 
32'd39280: dataIn1 = 32'd36
; 
32'd39281: dataIn1 = 32'd37
; 
32'd39282: dataIn1 = 32'd39
; 
32'd39283: dataIn1 = 32'd40
; 
32'd39284: dataIn1 = 32'd41
; 
32'd39285: dataIn1 = 32'd42
; 
32'd39286: dataIn1 = 32'd43
; 
32'd39287: dataIn1 = 32'd44
; 
32'd39288: dataIn1 = 32'd47
; 
32'd39289: dataIn1 = 32'd48
; 
32'd39290: dataIn1 = 32'd49
; 
32'd39291: dataIn1 = 32'd51
; 
32'd39292: dataIn1 = 32'd52
; 
32'd39293: dataIn1 = 32'd53
; 
32'd39294: dataIn1 = 32'd55
; 
32'd39295: dataIn1 = 32'd56
; 
32'd39296: dataIn1 = 32'd57
; 
32'd39297: dataIn1 = 32'd58
; 
32'd39298: dataIn1 = 32'd59
; 
32'd39299: dataIn1 = 32'd62
; 
32'd39300: dataIn1 = 32'd63
; 
32'd39301: dataIn1 = 32'd; 
32'd39302: dataIn1 = 32'd; 
32'd39303: dataIn1 = 32'd; 
32'd39304: dataIn1 = 32'd; 
32'd39305: dataIn1 = 32'd; 
32'd39306: dataIn1 = 32'd; 
32'd39307: dataIn1 = 32'd; 
32'd39308: dataIn1 = 32'd; 
32'd39309: dataIn1 = 32'd; 
32'd39310: dataIn1 = 32'd; 
32'd39311: dataIn1 = 32'd; 
32'd39312: dataIn1 = 32'd; 
32'd39313: dataIn1 = 32'd; 
32'd39314: dataIn1 = 32'd; 
32'd39315: dataIn1 = 32'd; 
32'd39316: dataIn1 = 32'd; 
32'd39317: dataIn1 = 32'd; 
32'd39318: dataIn1 = 32'd; 
32'd39319: dataIn1 = 32'd; 
32'd39320: dataIn1 = 32'd; 
32'd39321: dataIn1 = 32'd; 
32'd39322: dataIn1 = 32'd; 
32'd39323: dataIn1 = 32'd; 
32'd39324: dataIn1 = 32'd; 
32'd39325: dataIn1 = 32'd; 
32'd39326: dataIn1 = 32'd; 
32'd39327: dataIn1 = 32'd; 
32'd39328: dataIn1 = 32'd; 
32'd39329: dataIn1 = 32'd; 
32'd39330: dataIn1 = 32'd; 
32'd39331: dataIn1 = 32'd; 
32'd39332: dataIn1 = 32'd; 
32'd39333: dataIn1 = 32'd; 
32'd39334: dataIn1 = 32'd; 
32'd39335: dataIn1 = 32'd; 
32'd39336: dataIn1 = 32'd; 
32'd39337: dataIn1 = 32'd; 
32'd39338: dataIn1 = 32'd; 
32'd39339: dataIn1 = 32'd; 
32'd39340: dataIn1 = 32'd; 
32'd39341: dataIn1 = 32'd; 
32'd39342: dataIn1 = 32'd; 
32'd39343: dataIn1 = 32'd; 
32'd39344: dataIn1 = 32'd; 
32'd39345: dataIn1 = 32'd; 
32'd39346: dataIn1 = 32'd; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd23; 
32'd3: dataIn2 = 32'd62; 
32'd4: dataIn2 = 32'd2; 
32'd5: dataIn2 = 32'd39; 
32'd6: dataIn2 = 32'd93; 
32'd7: dataIn2 = 32'd19; 
32'd8: dataIn2 = 32'd31; 
32'd9: dataIn2 = 32'd15; 
32'd10: dataIn2 = 32'd48; 
32'd11: dataIn2 = 32'd50; 
32'd12: dataIn2 = 32'd0; 
32'd13: dataIn2 = 32'd26; 
32'd14: dataIn2 = 32'd87; 
32'd15: dataIn2 = 32'd89; 
32'd16: dataIn2 = 32'd96; 
32'd17: dataIn2 = 32'd57; 
32'd18: dataIn2 = 32'd18; 
32'd19: dataIn2 = 32'd71; 
32'd20: dataIn2 = 32'd75; 
32'd21: dataIn2 = 32'd79; 
32'd22: dataIn2 = 32'd0; 
32'd23: dataIn2 = 32'd82; 
32'd24: dataIn2 = 32'd2; 
32'd25: dataIn2 = 32'd65; 
32'd26: dataIn2 = 32'd40; 
32'd27: dataIn2 = 32'd78; 
32'd28: dataIn2 = 32'd0; 
32'd29: dataIn2 = 32'd77; 
32'd30: dataIn2 = 32'd42; 
32'd31: dataIn2 = 32'd44; 
32'd32: dataIn2 = 32'd74; 
32'd33: dataIn2 = 32'd93; 
32'd34: dataIn2 = 32'd83; 
32'd35: dataIn2 = 32'd4; 
32'd36: dataIn2 = 32'd13; 
32'd37: dataIn2 = 32'd61; 
32'd38: dataIn2 = 32'd59; 
32'd39: dataIn2 = 32'd47; 
32'd40: dataIn2 = 32'd20; 
32'd41: dataIn2 = 32'd84; 
32'd42: dataIn2 = 32'd17; 
32'd43: dataIn2 = 32'd70; 
32'd44: dataIn2 = 32'd69; 
32'd45: dataIn2 = 32'd90; 
32'd46: dataIn2 = 32'd46; 
32'd47: dataIn2 = 32'd59; 
32'd48: dataIn2 = 32'd76; 
32'd49: dataIn2 = 32'd1; 
32'd50: dataIn2 = 32'd28; 
32'd51: dataIn2 = 32'd54; 
32'd52: dataIn2 = 32'd23; 
32'd53: dataIn2 = 32'd10; 
32'd54: dataIn2 = 32'd27; 
32'd55: dataIn2 = 32'd33; 
32'd56: dataIn2 = 32'd52; 
32'd57: dataIn2 = 32'd22; 
32'd58: dataIn2 = 32'd16; 
32'd59: dataIn2 = 32'd25; 
32'd60: dataIn2 = 32'd90; 
32'd61: dataIn2 = 32'd10; 
32'd62: dataIn2 = 32'd28; 
32'd63: dataIn2 = 32'd59; 
32'd64: dataIn2 = 32'd68; 
32'd65: dataIn2 = 32'd15; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd330: dataIn2 = 32'd56; 
32'd331: dataIn2 = 32'd94; 
32'd332: dataIn2 = 32'd42; 
32'd333: dataIn2 = 32'd9; 
32'd334: dataIn2 = 32'd56; 
32'd335: dataIn2 = 32'd95; 
32'd336: dataIn2 = 32'd38; 
32'd337: dataIn2 = 32'd25; 
32'd338: dataIn2 = 32'd73; 
32'd339: dataIn2 = 32'd51; 
32'd340: dataIn2 = 32'd3; 
32'd341: dataIn2 = 32'd31; 
32'd342: dataIn2 = 32'd74; 
32'd343: dataIn2 = 32'd6; 
32'd344: dataIn2 = 32'd81; 
32'd345: dataIn2 = 32'd0; 
32'd346: dataIn2 = 32'd28; 
32'd347: dataIn2 = 32'd95; 
32'd348: dataIn2 = 32'd93; 
32'd349: dataIn2 = 32'd9; 
32'd350: dataIn2 = 32'd20; 
32'd351: dataIn2 = 32'd69; 
32'd352: dataIn2 = 32'd24; 
32'd353: dataIn2 = 32'd69; 
32'd354: dataIn2 = 32'd92; 
32'd355: dataIn2 = 32'd0; 
32'd356: dataIn2 = 32'd96; 
32'd357: dataIn2 = 32'd74; 
32'd358: dataIn2 = 32'd42; 
32'd359: dataIn2 = 32'd98; 
32'd360: dataIn2 = 32'd21; 
32'd361: dataIn2 = 32'd30; 
32'd362: dataIn2 = 32'd74; 
32'd363: dataIn2 = 32'd99; 
32'd364: dataIn2 = 32'd73; 
32'd365: dataIn2 = 32'd7; 
32'd366: dataIn2 = 32'd29; 
32'd367: dataIn2 = 32'd34; 
32'd368: dataIn2 = 32'd21; 
32'd369: dataIn2 = 32'd14; 
32'd370: dataIn2 = 32'd55; 
32'd371: dataIn2 = 32'd61; 
32'd372: dataIn2 = 32'd37; 
32'd373: dataIn2 = 32'd9; 
32'd374: dataIn2 = 32'd100; 
32'd375: dataIn2 = 32'd13; 
32'd376: dataIn2 = 32'd67; 
32'd377: dataIn2 = 32'd48; 
32'd378: dataIn2 = 32'd66; 
32'd379: dataIn2 = 32'd92; 
32'd380: dataIn2 = 32'd7; 
32'd381: dataIn2 = 32'd70; 
32'd382: dataIn2 = 32'd96; 
32'd383: dataIn2 = 32'd44; 
32'd384: dataIn2 = 32'd75; 
32'd385: dataIn2 = 32'd8; 
32'd386: dataIn2 = 32'd29; 
32'd387: dataIn2 = 32'd93; 
32'd388: dataIn2 = 32'd39; 
32'd389: dataIn2 = 32'd82; 
32'd390: dataIn2 = 32'd21; 
32'd391: dataIn2 = 32'd57; 
32'd392: dataIn2 = 32'd12; 
32'd393: dataIn2 = 32'd84; 
32'd394: dataIn2 = 32'd6; 
32'd395: dataIn2 = 32'd81; 
32'd396: dataIn2 = 32'd67; 
32'd397: dataIn2 = 32'd61; 
32'd398: dataIn2 = 32'd67; 
32'd399: dataIn2 = 32'd38; 
32'd400: dataIn2 = 32'd37; 
32'd401: dataIn2 = 32'd26; 
32'd402: dataIn2 = 32'd7; 
32'd403: dataIn2 = 32'd96; 
32'd404: dataIn2 = 32'd65; 
32'd405: dataIn2 = 32'd7; 
32'd406: dataIn2 = 32'd55; 
32'd407: dataIn2 = 32'd81; 
32'd408: dataIn2 = 32'd54; 
32'd409: dataIn2 = 32'd0; 
32'd410: dataIn2 = 32'd16; 
32'd411: dataIn2 = 32'd25; 
32'd412: dataIn2 = 32'd2; 
32'd413: dataIn2 = 32'd3; 
32'd414: dataIn2 = 32'd27; 
32'd415: dataIn2 = 32'd13; 
32'd416: dataIn2 = 32'd53; 
32'd417: dataIn2 = 32'd76; 
32'd418: dataIn2 = 32'd67; 
32'd419: dataIn2 = 32'd14; 
32'd420: dataIn2 = 32'd19; 
32'd421: dataIn2 = 32'd8; 
32'd422: dataIn2 = 32'd42; 
32'd423: dataIn2 = 32'd8; 
32'd424: dataIn2 = 32'd7; 
32'd425: dataIn2 = 32'd28; 
32'd426: dataIn2 = 32'd27; 
32'd427: dataIn2 = 32'd88; 
32'd428: dataIn2 = 32'd100; 
32'd429: dataIn2 = 32'd5; 
32'd430: dataIn2 = 32'd15; 
32'd431: dataIn2 = 32'd18; 
32'd432: dataIn2 = 32'd34; 
32'd433: dataIn2 = 32'd92; 
32'd434: dataIn2 = 32'd25; 
32'd435: dataIn2 = 32'd78; 
32'd436: dataIn2 = 32'd67; 
32'd437: dataIn2 = 32'd76; 
32'd438: dataIn2 = 32'd27; 
32'd439: dataIn2 = 32'd86; 
32'd440: dataIn2 = 32'd48; 
32'd441: dataIn2 = 32'd11; 
32'd442: dataIn2 = 32'd61; 
32'd443: dataIn2 = 32'd27; 
32'd444: dataIn2 = 32'd96; 
32'd445: dataIn2 = 32'd19; 
32'd446: dataIn2 = 32'd62; 
32'd447: dataIn2 = 32'd75; 
32'd448: dataIn2 = 32'd99; 
32'd449: dataIn2 = 32'd52; 
32'd450: dataIn2 = 32'd31; 
32'd451: dataIn2 = 32'd37; 
32'd452: dataIn2 = 32'd0; 
32'd453: dataIn2 = 32'd1; 
32'd454: dataIn2 = 32'd1; 
32'd455: dataIn2 = 32'd40; 
32'd456: dataIn2 = 32'd8; 
32'd457: dataIn2 = 32'd40; 
32'd458: dataIn2 = 32'd71; 
32'd459: dataIn2 = 32'd87; 
32'd460: dataIn2 = 32'd54; 
32'd461: dataIn2 = 32'd9; 
32'd462: dataIn2 = 32'd65; 
32'd463: dataIn2 = 32'd49; 
32'd464: dataIn2 = 32'd51; 
32'd465: dataIn2 = 32'd100; 
32'd466: dataIn2 = 32'd92; 
32'd467: dataIn2 = 32'd56; 
32'd468: dataIn2 = 32'd1; 
32'd469: dataIn2 = 32'd79; 
32'd470: dataIn2 = 32'd89; 
32'd471: dataIn2 = 32'd14; 
32'd472: dataIn2 = 32'd24; 
32'd473: dataIn2 = 32'd13; 
32'd474: dataIn2 = 32'd60; 
32'd475: dataIn2 = 32'd41; 
32'd476: dataIn2 = 32'd8; 
32'd477: dataIn2 = 32'd31; 
32'd478: dataIn2 = 32'd13; 
32'd479: dataIn2 = 32'd21; 
32'd480: dataIn2 = 32'd29; 
32'd481: dataIn2 = 32'd76; 
32'd482: dataIn2 = 32'd98; 
32'd483: dataIn2 = 32'd52; 
32'd484: dataIn2 = 32'd40; 
32'd485: dataIn2 = 32'd22; 
32'd486: dataIn2 = 32'd68; 
32'd487: dataIn2 = 32'd35; 
32'd488: dataIn2 = 32'd75; 
32'd489: dataIn2 = 32'd99; 
32'd490: dataIn2 = 32'd31; 
32'd491: dataIn2 = 32'd30; 
32'd492: dataIn2 = 32'd33; 
32'd493: dataIn2 = 32'd24; 
32'd494: dataIn2 = 32'd30; 
32'd495: dataIn2 = 32'd83; 
32'd496: dataIn2 = 32'd92; 
32'd497: dataIn2 = 32'd73; 
32'd498: dataIn2 = 32'd84; 
32'd499: dataIn2 = 32'd88; 
32'd500: dataIn2 = 32'd34; 
32'd501: dataIn2 = 32'd63; 
32'd502: dataIn2 = 32'd20; 
32'd503: dataIn2 = 32'd55; 
32'd504: dataIn2 = 32'd99; 
32'd505: dataIn2 = 32'd50; 
32'd506: dataIn2 = 32'd33; 
32'd507: dataIn2 = 32'd84; 
32'd508: dataIn2 = 32'd91; 
32'd509: dataIn2 = 32'd22; 
32'd510: dataIn2 = 32'd47; 
32'd511: dataIn2 = 32'd66; 
32'd512: dataIn2 = 32'd86; 
32'd513: dataIn2 = 32'd32; 
32'd514: dataIn2 = 32'd69; 
32'd515: dataIn2 = 32'd6; 
32'd516: dataIn2 = 32'd52; 
32'd517: dataIn2 = 32'd30; 
32'd518: dataIn2 = 32'd16; 
32'd519: dataIn2 = 32'd94; 
32'd520: dataIn2 = 32'd48; 
32'd521: dataIn2 = 32'd24; 
32'd522: dataIn2 = 32'd73; 
32'd523: dataIn2 = 32'd66; 
32'd524: dataIn2 = 32'd40; 
32'd525: dataIn2 = 32'd86; 
32'd526: dataIn2 = 32'd15; 
32'd527: dataIn2 = 32'd53; 
32'd528: dataIn2 = 32'd81; 
32'd529: dataIn2 = 32'd35; 
32'd530: dataIn2 = 32'd77; 
32'd531: dataIn2 = 32'd84; 
32'd532: dataIn2 = 32'd16; 
32'd533: dataIn2 = 32'd13; 
32'd534: dataIn2 = 32'd43; 
32'd535: dataIn2 = 32'd96; 
32'd536: dataIn2 = 32'd82; 
32'd537: dataIn2 = 32'd17; 
32'd538: dataIn2 = 32'd23; 
32'd539: dataIn2 = 32'd22; 
32'd540: dataIn2 = 32'd11; 
32'd541: dataIn2 = 32'd99; 
32'd542: dataIn2 = 32'd76; 
32'd543: dataIn2 = 32'd50; 
32'd544: dataIn2 = 32'd97; 
32'd545: dataIn2 = 32'd35; 
32'd546: dataIn2 = 32'd34; 
32'd547: dataIn2 = 32'd27; 
32'd548: dataIn2 = 32'd86; 
32'd549: dataIn2 = 32'd53; 
32'd550: dataIn2 = 32'd68; 
32'd551: dataIn2 = 32'd89; 
32'd552: dataIn2 = 32'd14; 
32'd553: dataIn2 = 32'd20; 
32'd554: dataIn2 = 32'd76; 
32'd555: dataIn2 = 32'd45; 
32'd556: dataIn2 = 32'd60; 
32'd557: dataIn2 = 32'd49; 
32'd558: dataIn2 = 32'd48; 
32'd559: dataIn2 = 32'd45; 
32'd560: dataIn2 = 32'd76; 
32'd561: dataIn2 = 32'd48; 
32'd562: dataIn2 = 32'd39; 
32'd563: dataIn2 = 32'd26; 
32'd564: dataIn2 = 32'd98; 
32'd565: dataIn2 = 32'd12; 
32'd566: dataIn2 = 32'd96; 
32'd567: dataIn2 = 32'd53; 
32'd568: dataIn2 = 32'd90; 
32'd569: dataIn2 = 32'd47; 
32'd570: dataIn2 = 32'd41; 
32'd571: dataIn2 = 32'd12; 
32'd572: dataIn2 = 32'd94; 
32'd573: dataIn2 = 32'd49; 
32'd574: dataIn2 = 32'd50; 
32'd575: dataIn2 = 32'd71; 
32'd576: dataIn2 = 32'd12; 
32'd577: dataIn2 = 32'd84; 
32'd578: dataIn2 = 32'd73; 
32'd579: dataIn2 = 32'd64; 
32'd580: dataIn2 = 32'd80; 
32'd581: dataIn2 = 32'd66; 
32'd582: dataIn2 = 32'd61; 
32'd583: dataIn2 = 32'd28; 
32'd584: dataIn2 = 32'd45; 
32'd585: dataIn2 = 32'd47; 
32'd586: dataIn2 = 32'd76; 
32'd587: dataIn2 = 32'd99; 
32'd588: dataIn2 = 32'd76; 
32'd589: dataIn2 = 32'd69; 
32'd590: dataIn2 = 32'd27; 
32'd591: dataIn2 = 32'd93; 
32'd592: dataIn2 = 32'd2; 
32'd593: dataIn2 = 32'd32; 
32'd594: dataIn2 = 32'd6; 
32'd595: dataIn2 = 32'd31; 
32'd596: dataIn2 = 32'd45; 
32'd597: dataIn2 = 32'd70; 
32'd598: dataIn2 = 32'd51; 
32'd599: dataIn2 = 32'd4; 
32'd600: dataIn2 = 32'd67; 
32'd601: dataIn2 = 32'd94; 
32'd602: dataIn2 = 32'd21; 
32'd603: dataIn2 = 32'd87; 
32'd604: dataIn2 = 32'd89; 
32'd605: dataIn2 = 32'd15; 
32'd606: dataIn2 = 32'd2; 
32'd607: dataIn2 = 32'd17; 
32'd608: dataIn2 = 32'd80; 
32'd609: dataIn2 = 32'd55; 
32'd610: dataIn2 = 32'd20; 
32'd611: dataIn2 = 32'd2; 
32'd612: dataIn2 = 32'd43; 
32'd613: dataIn2 = 32'd94; 
32'd614: dataIn2 = 32'd44; 
32'd615: dataIn2 = 32'd38; 
32'd616: dataIn2 = 32'd99; 
32'd617: dataIn2 = 32'd84; 
32'd618: dataIn2 = 32'd22; 
32'd619: dataIn2 = 32'd29; 
32'd620: dataIn2 = 32'd29; 
32'd621: dataIn2 = 32'd12; 
32'd622: dataIn2 = 32'd1; 
32'd623: dataIn2 = 32'd36; 
32'd624: dataIn2 = 32'd91; 
32'd625: dataIn2 = 32'd86; 
32'd626: dataIn2 = 32'd98; 
32'd627: dataIn2 = 32'd18; 
32'd628: dataIn2 = 32'd77; 
32'd629: dataIn2 = 32'd46; 
32'd630: dataIn2 = 32'd33; 
32'd631: dataIn2 = 32'd35; 
32'd632: dataIn2 = 32'd100; 
32'd633: dataIn2 = 32'd41; 
32'd634: dataIn2 = 32'd63; 
32'd635: dataIn2 = 32'd43; 
32'd636: dataIn2 = 32'd94; 
32'd637: dataIn2 = 32'd87; 
32'd638: dataIn2 = 32'd18; 
32'd639: dataIn2 = 32'd84; 
32'd640: dataIn2 = 32'd34; 
32'd641: dataIn2 = 32'd74; 
32'd642: dataIn2 = 32'd22; 
32'd643: dataIn2 = 32'd96; 
32'd644: dataIn2 = 32'd98; 
32'd645: dataIn2 = 32'd1; 
32'd646: dataIn2 = 32'd75; 
32'd647: dataIn2 = 32'd23; 
32'd648: dataIn2 = 32'd21; 
32'd649: dataIn2 = 32'd19; 
32'd650: dataIn2 = 32'd46; 
32'd651: dataIn2 = 32'd46; 
32'd652: dataIn2 = 32'd57; 
32'd653: dataIn2 = 32'd17; 
32'd654: dataIn2 = 32'd86; 
32'd655: dataIn2 = 32'd62; 
32'd656: dataIn2 = 32'd42; 
32'd657: dataIn2 = 32'd21; 
32'd658: dataIn2 = 32'd78; 
32'd659: dataIn2 = 32'd20; 
32'd660: dataIn2 = 32'd12; 
32'd661: dataIn2 = 32'd64; 
32'd662: dataIn2 = 32'd22; 
32'd663: dataIn2 = 32'd12; 
32'd664: dataIn2 = 32'd99; 
32'd665: dataIn2 = 32'd65; 
32'd666: dataIn2 = 32'd83; 
32'd667: dataIn2 = 32'd2; 
32'd668: dataIn2 = 32'd91; 
32'd669: dataIn2 = 32'd73; 
32'd670: dataIn2 = 32'd50; 
32'd671: dataIn2 = 32'd78; 
32'd672: dataIn2 = 32'd64; 
32'd673: dataIn2 = 32'd26; 
32'd674: dataIn2 = 32'd13; 
32'd675: dataIn2 = 32'd17; 
32'd676: dataIn2 = 32'd57; 
32'd677: dataIn2 = 32'd44; 
32'd678: dataIn2 = 32'd54; 
32'd679: dataIn2 = 32'd68; 
32'd680: dataIn2 = 32'd8; 
32'd681: dataIn2 = 32'd24; 
32'd682: dataIn2 = 32'd65; 
32'd683: dataIn2 = 32'd20; 
32'd684: dataIn2 = 32'd96; 
32'd685: dataIn2 = 32'd91; 
32'd686: dataIn2 = 32'd4; 
32'd687: dataIn2 = 32'd55; 
32'd688: dataIn2 = 32'd72; 
32'd689: dataIn2 = 32'd77; 
32'd690: dataIn2 = 32'd82; 
32'd691: dataIn2 = 32'd31; 
32'd692: dataIn2 = 32'd5; 
32'd693: dataIn2 = 32'd3; 
32'd694: dataIn2 = 32'd15; 
32'd695: dataIn2 = 32'd64; 
32'd696: dataIn2 = 32'd29; 
32'd697: dataIn2 = 32'd29; 
32'd698: dataIn2 = 32'd67; 
32'd699: dataIn2 = 32'd62; 
32'd700: dataIn2 = 32'd10; 
32'd701: dataIn2 = 32'd55; 
32'd702: dataIn2 = 32'd97; 
32'd703: dataIn2 = 32'd10; 
32'd704: dataIn2 = 32'd52; 
32'd705: dataIn2 = 32'd75; 
32'd706: dataIn2 = 32'd78; 
32'd707: dataIn2 = 32'd6; 
32'd708: dataIn2 = 32'd76; 
32'd709: dataIn2 = 32'd64; 
32'd710: dataIn2 = 32'd19; 
32'd711: dataIn2 = 32'd50; 
32'd712: dataIn2 = 32'd11; 
32'd713: dataIn2 = 32'd65; 
32'd714: dataIn2 = 32'd9; 
32'd715: dataIn2 = 32'd68; 
32'd716: dataIn2 = 32'd46; 
32'd717: dataIn2 = 32'd10; 
32'd718: dataIn2 = 32'd26; 
32'd719: dataIn2 = 32'd55; 
32'd720: dataIn2 = 32'd42; 
32'd721: dataIn2 = 32'd69; 
32'd722: dataIn2 = 32'd93; 
32'd723: dataIn2 = 32'd5; 
32'd724: dataIn2 = 32'd3; 
32'd725: dataIn2 = 32'd43; 
32'd726: dataIn2 = 32'd75; 
32'd727: dataIn2 = 32'd42; 
32'd728: dataIn2 = 32'd46; 
32'd729: dataIn2 = 32'd4; 
32'd730: dataIn2 = 32'd80; 
32'd731: dataIn2 = 32'd35; 
32'd732: dataIn2 = 32'd41; 
32'd733: dataIn2 = 32'd73; 
32'd734: dataIn2 = 32'd83; 
32'd735: dataIn2 = 32'd39; 
32'd736: dataIn2 = 32'd43; 
32'd737: dataIn2 = 32'd72; 
32'd738: dataIn2 = 32'd88; 
32'd739: dataIn2 = 32'd58; 
32'd740: dataIn2 = 32'd82; 
32'd741: dataIn2 = 32'd31; 
32'd742: dataIn2 = 32'd70; 
32'd743: dataIn2 = 32'd84; 
32'd744: dataIn2 = 32'd28; 
32'd745: dataIn2 = 32'd63; 
32'd746: dataIn2 = 32'd13; 
32'd747: dataIn2 = 32'd99; 
32'd748: dataIn2 = 32'd79; 
32'd749: dataIn2 = 32'd27; 
32'd750: dataIn2 = 32'd34; 
32'd751: dataIn2 = 32'd37; 
32'd752: dataIn2 = 32'd34; 
32'd753: dataIn2 = 32'd35; 
32'd754: dataIn2 = 32'd74; 
32'd755: dataIn2 = 32'd51; 
32'd756: dataIn2 = 32'd80; 
32'd757: dataIn2 = 32'd64; 
32'd758: dataIn2 = 32'd51; 
32'd759: dataIn2 = 32'd17; 
32'd760: dataIn2 = 32'd71; 
32'd761: dataIn2 = 32'd60; 
32'd762: dataIn2 = 32'd37; 
32'd763: dataIn2 = 32'd6; 
32'd764: dataIn2 = 32'd17; 
32'd765: dataIn2 = 32'd17; 
32'd766: dataIn2 = 32'd65; 
32'd767: dataIn2 = 32'd78; 
32'd768: dataIn2 = 32'd71; 
32'd769: dataIn2 = 32'd26; 
32'd770: dataIn2 = 32'd21; 
32'd771: dataIn2 = 32'd99; 
32'd772: dataIn2 = 32'd26; 
32'd773: dataIn2 = 32'd36; 
32'd774: dataIn2 = 32'd78; 
32'd775: dataIn2 = 32'd83; 
32'd776: dataIn2 = 32'd36; 
32'd777: dataIn2 = 32'd47; 
32'd778: dataIn2 = 32'd45; 
32'd779: dataIn2 = 32'd60; 
32'd780: dataIn2 = 32'd46; 
32'd781: dataIn2 = 32'd68; 
32'd782: dataIn2 = 32'd19; 
32'd783: dataIn2 = 32'd68; 
32'd784: dataIn2 = 32'd58; 
32'd785: dataIn2 = 32'd93; 
32'd786: dataIn2 = 32'd17; 
32'd787: dataIn2 = 32'd75; 
32'd788: dataIn2 = 32'd21; 
32'd789: dataIn2 = 32'd44; 
32'd790: dataIn2 = 32'd16; 
32'd791: dataIn2 = 32'd90; 
32'd792: dataIn2 = 32'd52; 
32'd793: dataIn2 = 32'd21; 
32'd794: dataIn2 = 32'd89; 
32'd795: dataIn2 = 32'd88; 
32'd796: dataIn2 = 32'd40; 
32'd797: dataIn2 = 32'd78; 
32'd798: dataIn2 = 32'd87; 
32'd799: dataIn2 = 32'd46; 
32'd800: dataIn2 = 32'd48; 
32'd801: dataIn2 = 32'd38; 
32'd802: dataIn2 = 32'd50; 
32'd803: dataIn2 = 32'd12; 
32'd804: dataIn2 = 32'd70; 
32'd805: dataIn2 = 32'd67; 
32'd806: dataIn2 = 32'd69; 
32'd807: dataIn2 = 32'd57; 
32'd808: dataIn2 = 32'd94; 
32'd809: dataIn2 = 32'd66; 
32'd810: dataIn2 = 32'd34; 
32'd811: dataIn2 = 32'd49; 
32'd812: dataIn2 = 32'd56; 
32'd813: dataIn2 = 32'd62; 
32'd814: dataIn2 = 32'd91; 
32'd815: dataIn2 = 32'd27; 
32'd816: dataIn2 = 32'd49; 
32'd817: dataIn2 = 32'd66; 
32'd818: dataIn2 = 32'd66; 
32'd819: dataIn2 = 32'd35; 
32'd820: dataIn2 = 32'd24; 
32'd821: dataIn2 = 32'd82; 
32'd822: dataIn2 = 32'd54; 
32'd823: dataIn2 = 32'd43; 
32'd824: dataIn2 = 32'd5; 
32'd825: dataIn2 = 32'd95; 
32'd826: dataIn2 = 32'd68; 
32'd827: dataIn2 = 32'd49; 
32'd828: dataIn2 = 32'd25; 
32'd829: dataIn2 = 32'd51; 
32'd830: dataIn2 = 32'd2; 
32'd831: dataIn2 = 32'd52; 
32'd832: dataIn2 = 32'd62; 
32'd833: dataIn2 = 32'd45; 
32'd834: dataIn2 = 32'd66; 
32'd835: dataIn2 = 32'd12; 
32'd836: dataIn2 = 32'd89; 
32'd837: dataIn2 = 32'd5; 
32'd838: dataIn2 = 32'd86; 
32'd839: dataIn2 = 32'd71; 
32'd840: dataIn2 = 32'd40; 
32'd841: dataIn2 = 32'd32; 
32'd842: dataIn2 = 32'd38; 
32'd843: dataIn2 = 32'd49; 
32'd844: dataIn2 = 32'd96; 
32'd845: dataIn2 = 32'd68; 
32'd846: dataIn2 = 32'd49; 
32'd847: dataIn2 = 32'd83; 
32'd848: dataIn2 = 32'd19; 
32'd849: dataIn2 = 32'd17; 
32'd850: dataIn2 = 32'd71; 
32'd851: dataIn2 = 32'd96; 
32'd852: dataIn2 = 32'd1; 
32'd853: dataIn2 = 32'd16; 
32'd854: dataIn2 = 32'd65; 
32'd855: dataIn2 = 32'd34; 
32'd856: dataIn2 = 32'd47; 
32'd857: dataIn2 = 32'd23; 
32'd858: dataIn2 = 32'd34; 
32'd859: dataIn2 = 32'd67; 
32'd860: dataIn2 = 32'd57; 
32'd861: dataIn2 = 32'd81; 
32'd862: dataIn2 = 32'd87; 
32'd863: dataIn2 = 32'd57; 
32'd864: dataIn2 = 32'd75; 
32'd865: dataIn2 = 32'd53; 
32'd866: dataIn2 = 32'd15; 
32'd867: dataIn2 = 32'd42; 
32'd868: dataIn2 = 32'd32; 
32'd869: dataIn2 = 32'd94; 
32'd870: dataIn2 = 32'd46; 
32'd871: dataIn2 = 32'd1; 
32'd872: dataIn2 = 32'd32; 
32'd873: dataIn2 = 32'd54; 
32'd874: dataIn2 = 32'd5; 
32'd875: dataIn2 = 32'd72; 
32'd876: dataIn2 = 32'd64; 
32'd877: dataIn2 = 32'd52; 
32'd878: dataIn2 = 32'd89; 
32'd879: dataIn2 = 32'd46; 
32'd880: dataIn2 = 32'd20; 
32'd881: dataIn2 = 32'd1; 
32'd882: dataIn2 = 32'd8; 
32'd883: dataIn2 = 32'd50; 
32'd884: dataIn2 = 32'd62; 
32'd885: dataIn2 = 32'd5; 
32'd886: dataIn2 = 32'd24; 
32'd887: dataIn2 = 32'd70; 
32'd888: dataIn2 = 32'd0; 
32'd889: dataIn2 = 32'd82; 
32'd890: dataIn2 = 32'd10; 
32'd891: dataIn2 = 32'd1; 
32'd892: dataIn2 = 32'd92; 
32'd893: dataIn2 = 32'd1; 
32'd894: dataIn2 = 32'd74; 
32'd895: dataIn2 = 32'd43; 
32'd896: dataIn2 = 32'd28; 
32'd897: dataIn2 = 32'd49; 
32'd898: dataIn2 = 32'd74; 
32'd899: dataIn2 = 32'd12; 
32'd900: dataIn2 = 32'd91; 
32'd901: dataIn2 = 32'd37; 
32'd902: dataIn2 = 32'd41; 
32'd903: dataIn2 = 32'd86; 
32'd904: dataIn2 = 32'd5; 
32'd905: dataIn2 = 32'd51; 
32'd906: dataIn2 = 32'd18; 
32'd907: dataIn2 = 32'd64; 
32'd908: dataIn2 = 32'd20; 
32'd909: dataIn2 = 32'd44; 
32'd910: dataIn2 = 32'd51; 
32'd911: dataIn2 = 32'd40; 
32'd912: dataIn2 = 32'd56; 
32'd913: dataIn2 = 32'd32; 
32'd914: dataIn2 = 32'd39; 
32'd915: dataIn2 = 32'd60; 
32'd916: dataIn2 = 32'd13; 
32'd917: dataIn2 = 32'd4; 
32'd918: dataIn2 = 32'd67; 
32'd919: dataIn2 = 32'd56; 
32'd920: dataIn2 = 32'd75; 
32'd921: dataIn2 = 32'd63; 
32'd922: dataIn2 = 32'd12; 
32'd923: dataIn2 = 32'd63; 
32'd924: dataIn2 = 32'd27; 
32'd925: dataIn2 = 32'd76; 
32'd926: dataIn2 = 32'd78; 
32'd927: dataIn2 = 32'd92; 
32'd928: dataIn2 = 32'd77; 
32'd929: dataIn2 = 32'd86; 
32'd930: dataIn2 = 32'd27; 
32'd931: dataIn2 = 32'd73; 
32'd932: dataIn2 = 32'd56; 
32'd933: dataIn2 = 32'd66; 
32'd934: dataIn2 = 32'd1; 
32'd935: dataIn2 = 32'd44; 
32'd936: dataIn2 = 32'd38; 
32'd937: dataIn2 = 32'd77; 
32'd938: dataIn2 = 32'd92; 
32'd939: dataIn2 = 32'd68; 
32'd940: dataIn2 = 32'd56; 
32'd941: dataIn2 = 32'd43; 
32'd942: dataIn2 = 32'd89; 
32'd943: dataIn2 = 32'd49; 
32'd944: dataIn2 = 32'd50; 
32'd945: dataIn2 = 32'd56; 
32'd946: dataIn2 = 32'd50; 
32'd947: dataIn2 = 32'd99; 
32'd948: dataIn2 = 32'd98; 
32'd949: dataIn2 = 32'd0; 
32'd950: dataIn2 = 32'd52; 
32'd951: dataIn2 = 32'd62; 
32'd952: dataIn2 = 32'd20; 
32'd953: dataIn2 = 32'd82; 
32'd954: dataIn2 = 32'd61; 
32'd955: dataIn2 = 32'd11; 
32'd956: dataIn2 = 32'd3; 
32'd957: dataIn2 = 32'd75; 
32'd958: dataIn2 = 32'd53; 
32'd959: dataIn2 = 32'd16; 
32'd960: dataIn2 = 32'd100; 
32'd961: dataIn2 = 32'd96; 
32'd962: dataIn2 = 32'd87; 
32'd963: dataIn2 = 32'd63; 
32'd964: dataIn2 = 32'd68; 
32'd965: dataIn2 = 32'd48; 
32'd966: dataIn2 = 32'd88; 
32'd967: dataIn2 = 32'd72; 
32'd968: dataIn2 = 32'd40; 
32'd969: dataIn2 = 32'd27; 
32'd970: dataIn2 = 32'd85; 
32'd971: dataIn2 = 32'd79; 
32'd972: dataIn2 = 32'd63; 
32'd973: dataIn2 = 32'd28; 
32'd974: dataIn2 = 32'd70; 
32'd975: dataIn2 = 32'd36; 
32'd976: dataIn2 = 32'd95; 
32'd977: dataIn2 = 32'd41; 
32'd978: dataIn2 = 32'd12; 
32'd979: dataIn2 = 32'd95; 
32'd980: dataIn2 = 32'd66; 
32'd981: dataIn2 = 32'd57; 
32'd982: dataIn2 = 32'd84; 
32'd983: dataIn2 = 32'd53; 
32'd984: dataIn2 = 32'd40; 
32'd985: dataIn2 = 32'd15; 
32'd986: dataIn2 = 32'd61; 
32'd987: dataIn2 = 32'd74; 
32'd988: dataIn2 = 32'd73; 
32'd989: dataIn2 = 32'd51; 
32'd990: dataIn2 = 32'd0; 
32'd991: dataIn2 = 32'd34; 
32'd992: dataIn2 = 32'd72; 
32'd993: dataIn2 = 32'd85; 
32'd994: dataIn2 = 32'd38; 
32'd995: dataIn2 = 32'd40; 
32'd996: dataIn2 = 32'd76; 
32'd997: dataIn2 = 32'd69; 
32'd998: dataIn2 = 32'd45; 
32'd999: dataIn2 = 32'd5; 
32'd1000: dataIn2 = 32'd28; 
32'd1001: dataIn2 = 32'd89; 
32'd1002: dataIn2 = 32'd35; 
32'd1003: dataIn2 = 32'd66; 
32'd1004: dataIn2 = 32'd66; 
32'd1005: dataIn2 = 32'd9; 
32'd1006: dataIn2 = 32'd90; 
32'd1007: dataIn2 = 32'd92; 
32'd1008: dataIn2 = 32'd20; 
32'd1009: dataIn2 = 32'd20; 
32'd1010: dataIn2 = 32'd79; 
32'd1011: dataIn2 = 32'd100; 
32'd1012: dataIn2 = 32'd59; 
32'd1013: dataIn2 = 32'd44; 
32'd1014: dataIn2 = 32'd34; 
32'd1015: dataIn2 = 32'd34; 
32'd1016: dataIn2 = 32'd59; 
32'd1017: dataIn2 = 32'd71; 
32'd1018: dataIn2 = 32'd41; 
32'd1019: dataIn2 = 32'd32; 
32'd1020: dataIn2 = 32'd31; 
32'd1021: dataIn2 = 32'd35; 
32'd1022: dataIn2 = 32'd82; 
32'd1023: dataIn2 = 32'd89; 
32'd1024: dataIn2 = 32'd24; 
32'd1025: dataIn2 = 32'd31; 
32'd1026: dataIn2 = 32'd9; 
32'd1027: dataIn2 = 32'd68; 
32'd1028: dataIn2 = 32'd76; 
32'd1029: dataIn2 = 32'd57; 
32'd1030: dataIn2 = 32'd1; 
32'd1031: dataIn2 = 32'd94; 
32'd1032: dataIn2 = 32'd100; 
32'd1033: dataIn2 = 32'd51; 
32'd1034: dataIn2 = 32'd34; 
32'd1035: dataIn2 = 32'd91; 
32'd1036: dataIn2 = 32'd49; 
32'd1037: dataIn2 = 32'd48; 
32'd1038: dataIn2 = 32'd54; 
32'd1039: dataIn2 = 32'd40; 
32'd1040: dataIn2 = 32'd20; 
32'd1041: dataIn2 = 32'd16; 
32'd1042: dataIn2 = 32'd47; 
32'd1043: dataIn2 = 32'd73; 
32'd1044: dataIn2 = 32'd21; 
32'd1045: dataIn2 = 32'd89; 
32'd1046: dataIn2 = 32'd73; 
32'd1047: dataIn2 = 32'd66; 
32'd1048: dataIn2 = 32'd65; 
32'd1049: dataIn2 = 32'd20; 
32'd1050: dataIn2 = 32'd93; 
32'd1051: dataIn2 = 32'd96; 
32'd1052: dataIn2 = 32'd84; 
32'd1053: dataIn2 = 32'd45; 
32'd1054: dataIn2 = 32'd9; 
32'd1055: dataIn2 = 32'd36; 
32'd1056: dataIn2 = 32'd16; 
32'd1057: dataIn2 = 32'd99; 
32'd1058: dataIn2 = 32'd30; 
32'd1059: dataIn2 = 32'd51; 
32'd1060: dataIn2 = 32'd98; 
32'd1061: dataIn2 = 32'd17; 
32'd1062: dataIn2 = 32'd91; 
32'd1063: dataIn2 = 32'd5; 
32'd1064: dataIn2 = 32'd79; 
32'd1065: dataIn2 = 32'd88; 
32'd1066: dataIn2 = 32'd52; 
32'd1067: dataIn2 = 32'd61; 
32'd1068: dataIn2 = 32'd64; 
32'd1069: dataIn2 = 32'd83; 
32'd1070: dataIn2 = 32'd32; 
32'd1071: dataIn2 = 32'd22; 
32'd1072: dataIn2 = 32'd92; 
32'd1073: dataIn2 = 32'd17; 
32'd1074: dataIn2 = 32'd23; 
32'd1075: dataIn2 = 32'd79; 
32'd1076: dataIn2 = 32'd63; 
32'd1077: dataIn2 = 32'd78; 
32'd1078: dataIn2 = 32'd72; 
32'd1079: dataIn2 = 32'd47; 
32'd1080: dataIn2 = 32'd89; 
32'd1081: dataIn2 = 32'd11; 
32'd1082: dataIn2 = 32'd17; 
32'd1083: dataIn2 = 32'd18; 
32'd1084: dataIn2 = 32'd85; 
32'd1085: dataIn2 = 32'd89; 
32'd1086: dataIn2 = 32'd87; 
32'd1087: dataIn2 = 32'd43; 
32'd1088: dataIn2 = 32'd2; 
32'd1089: dataIn2 = 32'd14; 
32'd1090: dataIn2 = 32'd87; 
32'd1091: dataIn2 = 32'd79; 
32'd1092: dataIn2 = 32'd64; 
32'd1093: dataIn2 = 32'd17; 
32'd1094: dataIn2 = 32'd53; 
32'd1095: dataIn2 = 32'd49; 
32'd1096: dataIn2 = 32'd81; 
32'd1097: dataIn2 = 32'd9; 
32'd1098: dataIn2 = 32'd76; 
32'd1099: dataIn2 = 32'd34; 
32'd1100: dataIn2 = 32'd57; 
32'd1101: dataIn2 = 32'd6; 
32'd1102: dataIn2 = 32'd45; 
32'd1103: dataIn2 = 32'd86; 
32'd1104: dataIn2 = 32'd51; 
32'd1105: dataIn2 = 32'd42; 
32'd1106: dataIn2 = 32'd60; 
32'd1107: dataIn2 = 32'd52; 
32'd1108: dataIn2 = 32'd35; 
32'd1109: dataIn2 = 32'd94; 
32'd1110: dataIn2 = 32'd98; 
32'd1111: dataIn2 = 32'd75; 
32'd1112: dataIn2 = 32'd57; 
32'd1113: dataIn2 = 32'd21; 
32'd1114: dataIn2 = 32'd83; 
32'd1115: dataIn2 = 32'd77; 
32'd1116: dataIn2 = 32'd77; 
32'd1117: dataIn2 = 32'd21; 
32'd1118: dataIn2 = 32'd32; 
32'd1119: dataIn2 = 32'd11; 
32'd1120: dataIn2 = 32'd48; 
32'd1121: dataIn2 = 32'd8; 
32'd1122: dataIn2 = 32'd27; 
32'd1123: dataIn2 = 32'd26; 
32'd1124: dataIn2 = 32'd40; 
32'd1125: dataIn2 = 32'd99; 
32'd1126: dataIn2 = 32'd89; 
32'd1127: dataIn2 = 32'd26; 
32'd1128: dataIn2 = 32'd66; 
32'd1129: dataIn2 = 32'd91; 
32'd1130: dataIn2 = 32'd26; 
32'd1131: dataIn2 = 32'd84; 
32'd1132: dataIn2 = 32'd58; 
32'd1133: dataIn2 = 32'd92; 
32'd1134: dataIn2 = 32'd50; 
32'd1135: dataIn2 = 32'd92; 
32'd1136: dataIn2 = 32'd93; 
32'd1137: dataIn2 = 32'd96; 
32'd1138: dataIn2 = 32'd29; 
32'd1139: dataIn2 = 32'd28; 
32'd1140: dataIn2 = 32'd37; 
32'd1141: dataIn2 = 32'd95; 
32'd1142: dataIn2 = 32'd20; 
32'd1143: dataIn2 = 32'd39; 
32'd1144: dataIn2 = 32'd24; 
32'd1145: dataIn2 = 32'd28; 
32'd1146: dataIn2 = 32'd28; 
32'd1147: dataIn2 = 32'd37; 
32'd1148: dataIn2 = 32'd18; 
32'd1149: dataIn2 = 32'd58; 
32'd1150: dataIn2 = 32'd47; 
32'd1151: dataIn2 = 32'd60; 
32'd1152: dataIn2 = 32'd70; 
32'd1153: dataIn2 = 32'd26; 
32'd1154: dataIn2 = 32'd72; 
32'd1155: dataIn2 = 32'd78; 
32'd1156: dataIn2 = 32'd48; 
32'd1157: dataIn2 = 32'd6; 
32'd1158: dataIn2 = 32'd93; 
32'd1159: dataIn2 = 32'd99; 
32'd1160: dataIn2 = 32'd40; 
32'd1161: dataIn2 = 32'd56; 
32'd1162: dataIn2 = 32'd59; 
32'd1163: dataIn2 = 32'd69; 
32'd1164: dataIn2 = 32'd54; 
32'd1165: dataIn2 = 32'd33; 
32'd1166: dataIn2 = 32'd16; 
32'd1167: dataIn2 = 32'd16; 
32'd1168: dataIn2 = 32'd23; 
32'd1169: dataIn2 = 32'd49; 
32'd1170: dataIn2 = 32'd25; 
32'd1171: dataIn2 = 32'd5; 
32'd1172: dataIn2 = 32'd40; 
32'd1173: dataIn2 = 32'd87; 
32'd1174: dataIn2 = 32'd48; 
32'd1175: dataIn2 = 32'd0; 
32'd1176: dataIn2 = 32'd69; 
32'd1177: dataIn2 = 32'd74; 
32'd1178: dataIn2 = 32'd81; 
32'd1179: dataIn2 = 32'd75; 
32'd1180: dataIn2 = 32'd94; 
32'd1181: dataIn2 = 32'd19; 
32'd1182: dataIn2 = 32'd54; 
32'd1183: dataIn2 = 32'd45; 
32'd1184: dataIn2 = 32'd73; 
32'd1185: dataIn2 = 32'd39; 
32'd1186: dataIn2 = 32'd77; 
32'd1187: dataIn2 = 32'd54; 
32'd1188: dataIn2 = 32'd30; 
32'd1189: dataIn2 = 32'd40; 
32'd1190: dataIn2 = 32'd19; 
32'd1191: dataIn2 = 32'd56; 
32'd1192: dataIn2 = 32'd55; 
32'd1193: dataIn2 = 32'd10; 
32'd1194: dataIn2 = 32'd77; 
32'd1195: dataIn2 = 32'd15; 
32'd1196: dataIn2 = 32'd16; 
32'd1197: dataIn2 = 32'd89; 
32'd1198: dataIn2 = 32'd33; 
32'd1199: dataIn2 = 32'd20; 
32'd1200: dataIn2 = 32'd76; 
32'd1201: dataIn2 = 32'd25; 
32'd1202: dataIn2 = 32'd87; 
32'd1203: dataIn2 = 32'd5; 
32'd1204: dataIn2 = 32'd45; 
32'd1205: dataIn2 = 32'd85; 
32'd1206: dataIn2 = 32'd65; 
32'd1207: dataIn2 = 32'd91; 
32'd1208: dataIn2 = 32'd85; 
32'd1209: dataIn2 = 32'd89; 
32'd1210: dataIn2 = 32'd8; 
32'd1211: dataIn2 = 32'd35; 
32'd1212: dataIn2 = 32'd86; 
32'd1213: dataIn2 = 32'd66; 
32'd1214: dataIn2 = 32'd83; 
32'd1215: dataIn2 = 32'd22; 
32'd1216: dataIn2 = 32'd68; 
32'd1217: dataIn2 = 32'd94; 
32'd1218: dataIn2 = 32'd21; 
32'd1219: dataIn2 = 32'd4; 
32'd1220: dataIn2 = 32'd18; 
32'd1221: dataIn2 = 32'd9; 
32'd1222: dataIn2 = 32'd49; 
32'd1223: dataIn2 = 32'd5; 
32'd1224: dataIn2 = 32'd42; 
32'd1225: dataIn2 = 32'd50; 
32'd1226: dataIn2 = 32'd61; 
32'd1227: dataIn2 = 32'd86; 
32'd1228: dataIn2 = 32'd47; 
32'd1229: dataIn2 = 32'd68; 
32'd1230: dataIn2 = 32'd58; 
32'd1231: dataIn2 = 32'd54; 
32'd1232: dataIn2 = 32'd93; 
32'd1233: dataIn2 = 32'd27; 
32'd1234: dataIn2 = 32'd77; 
32'd1235: dataIn2 = 32'd59; 
32'd1236: dataIn2 = 32'd2; 
32'd1237: dataIn2 = 32'd74; 
32'd1238: dataIn2 = 32'd29; 
32'd1239: dataIn2 = 32'd47; 
32'd1240: dataIn2 = 32'd23; 
32'd1241: dataIn2 = 32'd82; 
32'd1242: dataIn2 = 32'd52; 
32'd1243: dataIn2 = 32'd95; 
32'd1244: dataIn2 = 32'd74; 
32'd1245: dataIn2 = 32'd96; 
32'd1246: dataIn2 = 32'd61; 
32'd1247: dataIn2 = 32'd29; 
32'd1248: dataIn2 = 32'd97; 
32'd1249: dataIn2 = 32'd28; 
32'd1250: dataIn2 = 32'd58; 
32'd1251: dataIn2 = 32'd5; 
32'd1252: dataIn2 = 32'd29; 
32'd1253: dataIn2 = 32'd34; 
32'd1254: dataIn2 = 32'd92; 
32'd1255: dataIn2 = 32'd77; 
32'd1256: dataIn2 = 32'd94; 
32'd1257: dataIn2 = 32'd69; 
32'd1258: dataIn2 = 32'd3; 
32'd1259: dataIn2 = 32'd2; 
32'd1260: dataIn2 = 32'd2; 
32'd1261: dataIn2 = 32'd97; 
32'd1262: dataIn2 = 32'd48; 
32'd1263: dataIn2 = 32'd31; 
32'd1264: dataIn2 = 32'd37; 
32'd1265: dataIn2 = 32'd58; 
32'd1266: dataIn2 = 32'd98; 
32'd1267: dataIn2 = 32'd94; 
32'd1268: dataIn2 = 32'd71; 
32'd1269: dataIn2 = 32'd12; 
32'd1270: dataIn2 = 32'd37; 
32'd1271: dataIn2 = 32'd5; 
32'd1272: dataIn2 = 32'd83; 
32'd1273: dataIn2 = 32'd0; 
32'd1274: dataIn2 = 32'd68; 
32'd1275: dataIn2 = 32'd5; 
32'd1276: dataIn2 = 32'd22; 
32'd1277: dataIn2 = 32'd55; 
32'd1278: dataIn2 = 32'd57; 
32'd1279: dataIn2 = 32'd91; 
32'd1280: dataIn2 = 32'd25; 
32'd1281: dataIn2 = 32'd83; 
32'd1282: dataIn2 = 32'd5; 
32'd1283: dataIn2 = 32'd44; 
32'd1284: dataIn2 = 32'd13; 
32'd1285: dataIn2 = 32'd75; 
32'd1286: dataIn2 = 32'd8; 
32'd1287: dataIn2 = 32'd88; 
32'd1288: dataIn2 = 32'd26; 
32'd1289: dataIn2 = 32'd28; 
32'd1290: dataIn2 = 32'd8; 
32'd1291: dataIn2 = 32'd30; 
32'd1292: dataIn2 = 32'd77; 
32'd1293: dataIn2 = 32'd67; 
32'd1294: dataIn2 = 32'd14; 
32'd1295: dataIn2 = 32'd55; 
32'd1296: dataIn2 = 32'd45; 
32'd1297: dataIn2 = 32'd45; 
32'd1298: dataIn2 = 32'd78; 
32'd1299: dataIn2 = 32'd38; 
32'd1300: dataIn2 = 32'd28; 
32'd1301: dataIn2 = 32'd58; 
32'd1302: dataIn2 = 32'd0; 
32'd1303: dataIn2 = 32'd18; 
32'd1304: dataIn2 = 32'd85; 
32'd1305: dataIn2 = 32'd95; 
32'd1306: dataIn2 = 32'd51; 
32'd1307: dataIn2 = 32'd25; 
32'd1308: dataIn2 = 32'd4; 
32'd1309: dataIn2 = 32'd89; 
32'd1310: dataIn2 = 32'd77; 
32'd1311: dataIn2 = 32'd15; 
32'd1312: dataIn2 = 32'd60; 
32'd1313: dataIn2 = 32'd41; 
32'd1314: dataIn2 = 32'd94; 
32'd1315: dataIn2 = 32'd70; 
32'd1316: dataIn2 = 32'd66; 
32'd1317: dataIn2 = 32'd96; 
32'd1318: dataIn2 = 32'd49; 
32'd1319: dataIn2 = 32'd79; 
32'd1320: dataIn2 = 32'd85; 
32'd1321: dataIn2 = 32'd21; 
32'd1322: dataIn2 = 32'd49; 
32'd1323: dataIn2 = 32'd16; 
32'd1324: dataIn2 = 32'd5; 
32'd1325: dataIn2 = 32'd39; 
32'd1326: dataIn2 = 32'd34; 
32'd1327: dataIn2 = 32'd45; 
32'd1328: dataIn2 = 32'd35; 
32'd1329: dataIn2 = 32'd95; 
32'd1330: dataIn2 = 32'd34; 
32'd1331: dataIn2 = 32'd30; 
32'd1332: dataIn2 = 32'd10; 
32'd1333: dataIn2 = 32'd75; 
32'd1334: dataIn2 = 32'd5; 
32'd1335: dataIn2 = 32'd26; 
32'd1336: dataIn2 = 32'd35; 
32'd1337: dataIn2 = 32'd47; 
32'd1338: dataIn2 = 32'd73; 
32'd1339: dataIn2 = 32'd86; 
32'd1340: dataIn2 = 32'd29; 
32'd1341: dataIn2 = 32'd11; 
32'd1342: dataIn2 = 32'd10; 
32'd1343: dataIn2 = 32'd4; 
32'd1344: dataIn2 = 32'd14; 
32'd1345: dataIn2 = 32'd90; 
32'd1346: dataIn2 = 32'd3; 
32'd1347: dataIn2 = 32'd44; 
32'd1348: dataIn2 = 32'd6; 
32'd1349: dataIn2 = 32'd53; 
32'd1350: dataIn2 = 32'd30; 
32'd1351: dataIn2 = 32'd91; 
32'd1352: dataIn2 = 32'd38; 
32'd1353: dataIn2 = 32'd99; 
32'd1354: dataIn2 = 32'd87; 
32'd1355: dataIn2 = 32'd75; 
32'd1356: dataIn2 = 32'd23; 
32'd1357: dataIn2 = 32'd10; 
32'd1358: dataIn2 = 32'd5; 
32'd1359: dataIn2 = 32'd61; 
32'd1360: dataIn2 = 32'd96; 
32'd1361: dataIn2 = 32'd48; 
32'd1362: dataIn2 = 32'd46; 
32'd1363: dataIn2 = 32'd21; 
32'd1364: dataIn2 = 32'd72; 
32'd1365: dataIn2 = 32'd96; 
32'd1366: dataIn2 = 32'd83; 
32'd1367: dataIn2 = 32'd37; 
32'd1368: dataIn2 = 32'd64; 
32'd1369: dataIn2 = 32'd6; 
32'd1370: dataIn2 = 32'd51; 
32'd1371: dataIn2 = 32'd9; 
32'd1372: dataIn2 = 32'd38; 
32'd1373: dataIn2 = 32'd96; 
32'd1374: dataIn2 = 32'd47; 
32'd1375: dataIn2 = 32'd58; 
32'd1376: dataIn2 = 32'd33; 
32'd1377: dataIn2 = 32'd36; 
32'd1378: dataIn2 = 32'd10; 
32'd1379: dataIn2 = 32'd63; 
32'd1380: dataIn2 = 32'd10; 
32'd1381: dataIn2 = 32'd95; 
32'd1382: dataIn2 = 32'd82; 
32'd1383: dataIn2 = 32'd35; 
32'd1384: dataIn2 = 32'd12; 
32'd1385: dataIn2 = 32'd41; 
32'd1386: dataIn2 = 32'd81; 
32'd1387: dataIn2 = 32'd53; 
32'd1388: dataIn2 = 32'd77; 
32'd1389: dataIn2 = 32'd52; 
32'd1390: dataIn2 = 32'd89; 
32'd1391: dataIn2 = 32'd48; 
32'd1392: dataIn2 = 32'd96; 
32'd1393: dataIn2 = 32'd89; 
32'd1394: dataIn2 = 32'd67; 
32'd1395: dataIn2 = 32'd5; 
32'd1396: dataIn2 = 32'd97; 
32'd1397: dataIn2 = 32'd89; 
32'd1398: dataIn2 = 32'd62; 
32'd1399: dataIn2 = 32'd68; 
32'd1400: dataIn2 = 32'd10; 
32'd1401: dataIn2 = 32'd35; 
32'd1402: dataIn2 = 32'd48; 
32'd1403: dataIn2 = 32'd38; 
32'd1404: dataIn2 = 32'd62; 
32'd1405: dataIn2 = 32'd90; 
32'd1406: dataIn2 = 32'd90; 
32'd1407: dataIn2 = 32'd70; 
32'd1408: dataIn2 = 32'd5; 
32'd1409: dataIn2 = 32'd15; 
32'd1410: dataIn2 = 32'd26; 
32'd1411: dataIn2 = 32'd92; 
32'd1412: dataIn2 = 32'd8; 
32'd1413: dataIn2 = 32'd25; 
32'd1414: dataIn2 = 32'd57; 
32'd1415: dataIn2 = 32'd60; 
32'd1416: dataIn2 = 32'd32; 
32'd1417: dataIn2 = 32'd54; 
32'd1418: dataIn2 = 32'd49; 
32'd1419: dataIn2 = 32'd47; 
32'd1420: dataIn2 = 32'd23; 
32'd1421: dataIn2 = 32'd90; 
32'd1422: dataIn2 = 32'd1; 
32'd1423: dataIn2 = 32'd86; 
32'd1424: dataIn2 = 32'd62; 
32'd1425: dataIn2 = 32'd42; 
32'd1426: dataIn2 = 32'd32; 
32'd1427: dataIn2 = 32'd87; 
32'd1428: dataIn2 = 32'd1; 
32'd1429: dataIn2 = 32'd49; 
32'd1430: dataIn2 = 32'd96; 
32'd1431: dataIn2 = 32'd48; 
32'd1432: dataIn2 = 32'd6; 
32'd1433: dataIn2 = 32'd44; 
32'd1434: dataIn2 = 32'd78; 
32'd1435: dataIn2 = 32'd82; 
32'd1436: dataIn2 = 32'd21; 
32'd1437: dataIn2 = 32'd83; 
32'd1438: dataIn2 = 32'd18; 
32'd1439: dataIn2 = 32'd36; 
32'd1440: dataIn2 = 32'd0; 
32'd1441: dataIn2 = 32'd72; 
32'd1442: dataIn2 = 32'd30; 
32'd1443: dataIn2 = 32'd86; 
32'd1444: dataIn2 = 32'd9; 
32'd1445: dataIn2 = 32'd73; 
32'd1446: dataIn2 = 32'd54; 
32'd1447: dataIn2 = 32'd10; 
32'd1448: dataIn2 = 32'd89; 
32'd1449: dataIn2 = 32'd26; 
32'd1450: dataIn2 = 32'd66; 
32'd1451: dataIn2 = 32'd35; 
32'd1452: dataIn2 = 32'd0; 
32'd1453: dataIn2 = 32'd25; 
32'd1454: dataIn2 = 32'd31; 
32'd1455: dataIn2 = 32'd39; 
32'd1456: dataIn2 = 32'd97; 
32'd1457: dataIn2 = 32'd80; 
32'd1458: dataIn2 = 32'd31; 
32'd1459: dataIn2 = 32'd13; 
32'd1460: dataIn2 = 32'd44; 
32'd1461: dataIn2 = 32'd29; 
32'd1462: dataIn2 = 32'd46; 
32'd1463: dataIn2 = 32'd71; 
32'd1464: dataIn2 = 32'd91; 
32'd1465: dataIn2 = 32'd64; 
32'd1466: dataIn2 = 32'd74; 
32'd1467: dataIn2 = 32'd50; 
32'd1468: dataIn2 = 32'd18; 
32'd1469: dataIn2 = 32'd61; 
32'd1470: dataIn2 = 32'd97; 
32'd1471: dataIn2 = 32'd13; 
32'd1472: dataIn2 = 32'd35; 
32'd1473: dataIn2 = 32'd14; 
32'd1474: dataIn2 = 32'd13; 
32'd1475: dataIn2 = 32'd91; 
32'd1476: dataIn2 = 32'd29; 
32'd1477: dataIn2 = 32'd66; 
32'd1478: dataIn2 = 32'd2; 
32'd1479: dataIn2 = 32'd100; 
32'd1480: dataIn2 = 32'd69; 
32'd1481: dataIn2 = 32'd27; 
32'd1482: dataIn2 = 32'd100; 
32'd1483: dataIn2 = 32'd97; 
32'd1484: dataIn2 = 32'd52; 
32'd1485: dataIn2 = 32'd96; 
32'd1486: dataIn2 = 32'd14; 
32'd1487: dataIn2 = 32'd64; 
32'd1488: dataIn2 = 32'd99; 
32'd1489: dataIn2 = 32'd97; 
32'd1490: dataIn2 = 32'd56; 
32'd1491: dataIn2 = 32'd14; 
32'd1492: dataIn2 = 32'd72; 
32'd1493: dataIn2 = 32'd7; 
32'd1494: dataIn2 = 32'd85; 
32'd1495: dataIn2 = 32'd58; 
32'd1496: dataIn2 = 32'd10; 
32'd1497: dataIn2 = 32'd83; 
32'd1498: dataIn2 = 32'd94; 
32'd1499: dataIn2 = 32'd16; 
32'd1500: dataIn2 = 32'd13; 
32'd1501: dataIn2 = 32'd83; 
32'd1502: dataIn2 = 32'd34; 
32'd1503: dataIn2 = 32'd32; 
32'd1504: dataIn2 = 32'd90; 
32'd1505: dataIn2 = 32'd8; 
32'd1506: dataIn2 = 32'd25; 
32'd1507: dataIn2 = 32'd36; 
32'd1508: dataIn2 = 32'd33; 
32'd1509: dataIn2 = 32'd75; 
32'd1510: dataIn2 = 32'd21; 
32'd1511: dataIn2 = 32'd29; 
32'd1512: dataIn2 = 32'd44; 
32'd1513: dataIn2 = 32'd90; 
32'd1514: dataIn2 = 32'd11; 
32'd1515: dataIn2 = 32'd43; 
32'd1516: dataIn2 = 32'd30; 
32'd1517: dataIn2 = 32'd10; 
32'd1518: dataIn2 = 32'd100; 
32'd1519: dataIn2 = 32'd5; 
32'd1520: dataIn2 = 32'd52; 
32'd1521: dataIn2 = 32'd66; 
32'd1522: dataIn2 = 32'd61; 
32'd1523: dataIn2 = 32'd74; 
32'd1524: dataIn2 = 32'd45; 
32'd1525: dataIn2 = 32'd75; 
32'd1526: dataIn2 = 32'd19; 
32'd1527: dataIn2 = 32'd12; 
32'd1528: dataIn2 = 32'd42; 
32'd1529: dataIn2 = 32'd36; 
32'd1530: dataIn2 = 32'd43; 
32'd1531: dataIn2 = 32'd64; 
32'd1532: dataIn2 = 32'd93; 
32'd1533: dataIn2 = 32'd12; 
32'd1534: dataIn2 = 32'd19; 
32'd1535: dataIn2 = 32'd9; 
32'd1536: dataIn2 = 32'd41; 
32'd1537: dataIn2 = 32'd56; 
32'd1538: dataIn2 = 32'd8; 
32'd1539: dataIn2 = 32'd74; 
32'd1540: dataIn2 = 32'd69; 
32'd1541: dataIn2 = 32'd12; 
32'd1542: dataIn2 = 32'd74; 
32'd1543: dataIn2 = 32'd71; 
32'd1544: dataIn2 = 32'd31; 
32'd1545: dataIn2 = 32'd36; 
32'd1546: dataIn2 = 32'd37; 
32'd1547: dataIn2 = 32'd45; 
32'd1548: dataIn2 = 32'd72; 
32'd1549: dataIn2 = 32'd25; 
32'd1550: dataIn2 = 32'd7; 
32'd1551: dataIn2 = 32'd37; 
32'd1552: dataIn2 = 32'd83; 
32'd1553: dataIn2 = 32'd40; 
32'd1554: dataIn2 = 32'd95; 
32'd1555: dataIn2 = 32'd3; 
32'd1556: dataIn2 = 32'd0; 
32'd1557: dataIn2 = 32'd69; 
32'd1558: dataIn2 = 32'd11; 
32'd1559: dataIn2 = 32'd20; 
32'd1560: dataIn2 = 32'd87; 
32'd1561: dataIn2 = 32'd9; 
32'd1562: dataIn2 = 32'd68; 
32'd1563: dataIn2 = 32'd68; 
32'd1564: dataIn2 = 32'd27; 
32'd1565: dataIn2 = 32'd15; 
32'd1566: dataIn2 = 32'd34; 
32'd1567: dataIn2 = 32'd33; 
32'd1568: dataIn2 = 32'd89; 
32'd1569: dataIn2 = 32'd98; 
32'd1570: dataIn2 = 32'd0; 
32'd1571: dataIn2 = 32'd41; 
32'd1572: dataIn2 = 32'd35; 
32'd1573: dataIn2 = 32'd94; 
32'd1574: dataIn2 = 32'd75; 
32'd1575: dataIn2 = 32'd56; 
32'd1576: dataIn2 = 32'd26; 
32'd1577: dataIn2 = 32'd39; 
32'd1578: dataIn2 = 32'd33; 
32'd1579: dataIn2 = 32'd36; 
32'd1580: dataIn2 = 32'd69; 
32'd1581: dataIn2 = 32'd57; 
32'd1582: dataIn2 = 32'd1; 
32'd1583: dataIn2 = 32'd29; 
32'd1584: dataIn2 = 32'd62; 
32'd1585: dataIn2 = 32'd48; 
32'd1586: dataIn2 = 32'd40; 
32'd1587: dataIn2 = 32'd84; 
32'd1588: dataIn2 = 32'd46; 
32'd1589: dataIn2 = 32'd29; 
32'd1590: dataIn2 = 32'd29; 
32'd1591: dataIn2 = 32'd24; 
32'd1592: dataIn2 = 32'd82; 
32'd1593: dataIn2 = 32'd24; 
32'd1594: dataIn2 = 32'd72; 
32'd1595: dataIn2 = 32'd75; 
32'd1596: dataIn2 = 32'd39; 
32'd1597: dataIn2 = 32'd87; 
32'd1598: dataIn2 = 32'd55; 
32'd1599: dataIn2 = 32'd44; 
32'd1600: dataIn2 = 32'd25; 
32'd1601: dataIn2 = 32'd69; 
32'd1602: dataIn2 = 32'd75; 
32'd1603: dataIn2 = 32'd26; 
32'd1604: dataIn2 = 32'd45; 
32'd1605: dataIn2 = 32'd52; 
32'd1606: dataIn2 = 32'd50; 
32'd1607: dataIn2 = 32'd45; 
32'd1608: dataIn2 = 32'd18; 
32'd1609: dataIn2 = 32'd94; 
32'd1610: dataIn2 = 32'd93; 
32'd1611: dataIn2 = 32'd62; 
32'd1612: dataIn2 = 32'd41; 
32'd1613: dataIn2 = 32'd25; 
32'd1614: dataIn2 = 32'd24; 
32'd1615: dataIn2 = 32'd89; 
32'd1616: dataIn2 = 32'd39; 
32'd1617: dataIn2 = 32'd37; 
32'd1618: dataIn2 = 32'd46; 
32'd1619: dataIn2 = 32'd100; 
32'd1620: dataIn2 = 32'd42; 
32'd1621: dataIn2 = 32'd91; 
32'd1622: dataIn2 = 32'd57; 
32'd1623: dataIn2 = 32'd71; 
32'd1624: dataIn2 = 32'd36; 
32'd1625: dataIn2 = 32'd69; 
32'd1626: dataIn2 = 32'd100; 
32'd1627: dataIn2 = 32'd22; 
32'd1628: dataIn2 = 32'd64; 
32'd1629: dataIn2 = 32'd92; 
32'd1630: dataIn2 = 32'd28; 
32'd1631: dataIn2 = 32'd14; 
32'd1632: dataIn2 = 32'd23; 
32'd1633: dataIn2 = 32'd32; 
32'd1634: dataIn2 = 32'd48; 
32'd1635: dataIn2 = 32'd0; 
32'd1636: dataIn2 = 32'd31; 
32'd1637: dataIn2 = 32'd29; 
32'd1638: dataIn2 = 32'd70; 
32'd1639: dataIn2 = 32'd40; 
32'd1640: dataIn2 = 32'd16; 
32'd1641: dataIn2 = 32'd87; 
32'd1642: dataIn2 = 32'd31; 
32'd1643: dataIn2 = 32'd95; 
32'd1644: dataIn2 = 32'd19; 
32'd1645: dataIn2 = 32'd47; 
32'd1646: dataIn2 = 32'd19; 
32'd1647: dataIn2 = 32'd81; 
32'd1648: dataIn2 = 32'd71; 
32'd1649: dataIn2 = 32'd55; 
32'd1650: dataIn2 = 32'd33; 
32'd1651: dataIn2 = 32'd87; 
32'd1652: dataIn2 = 32'd33; 
32'd1653: dataIn2 = 32'd99; 
32'd1654: dataIn2 = 32'd13; 
32'd1655: dataIn2 = 32'd47; 
32'd1656: dataIn2 = 32'd75; 
32'd1657: dataIn2 = 32'd49; 
32'd1658: dataIn2 = 32'd100; 
32'd1659: dataIn2 = 32'd95; 
32'd1660: dataIn2 = 32'd17; 
32'd1661: dataIn2 = 32'd42; 
32'd1662: dataIn2 = 32'd25; 
32'd1663: dataIn2 = 32'd88; 
32'd1664: dataIn2 = 32'd24; 
32'd1665: dataIn2 = 32'd76; 
32'd1666: dataIn2 = 32'd50; 
32'd1667: dataIn2 = 32'd91; 
32'd1668: dataIn2 = 32'd16; 
32'd1669: dataIn2 = 32'd78; 
32'd1670: dataIn2 = 32'd38; 
32'd1671: dataIn2 = 32'd85; 
32'd1672: dataIn2 = 32'd63; 
32'd1673: dataIn2 = 32'd29; 
32'd1674: dataIn2 = 32'd33; 
32'd1675: dataIn2 = 32'd32; 
32'd1676: dataIn2 = 32'd31; 
32'd1677: dataIn2 = 32'd97; 
32'd1678: dataIn2 = 32'd72; 
32'd1679: dataIn2 = 32'd69; 
32'd1680: dataIn2 = 32'd42; 
32'd1681: dataIn2 = 32'd35; 
32'd1682: dataIn2 = 32'd61; 
32'd1683: dataIn2 = 32'd40; 
32'd1684: dataIn2 = 32'd83; 
32'd1685: dataIn2 = 32'd32; 
32'd1686: dataIn2 = 32'd59; 
32'd1687: dataIn2 = 32'd74; 
32'd1688: dataIn2 = 32'd53; 
32'd1689: dataIn2 = 32'd65; 
32'd1690: dataIn2 = 32'd77; 
32'd1691: dataIn2 = 32'd94; 
32'd1692: dataIn2 = 32'd42; 
32'd1693: dataIn2 = 32'd68; 
32'd1694: dataIn2 = 32'd39; 
32'd1695: dataIn2 = 32'd72; 
32'd1696: dataIn2 = 32'd79; 
32'd1697: dataIn2 = 32'd76; 
32'd1698: dataIn2 = 32'd39; 
32'd1699: dataIn2 = 32'd52; 
32'd1700: dataIn2 = 32'd10; 
32'd1701: dataIn2 = 32'd14; 
32'd1702: dataIn2 = 32'd56; 
32'd1703: dataIn2 = 32'd88; 
32'd1704: dataIn2 = 32'd75; 
32'd1705: dataIn2 = 32'd92; 
32'd1706: dataIn2 = 32'd35; 
32'd1707: dataIn2 = 32'd100; 
32'd1708: dataIn2 = 32'd57; 
32'd1709: dataIn2 = 32'd57; 
32'd1710: dataIn2 = 32'd34; 
32'd1711: dataIn2 = 32'd91; 
32'd1712: dataIn2 = 32'd17; 
32'd1713: dataIn2 = 32'd13; 
32'd1714: dataIn2 = 32'd16; 
32'd1715: dataIn2 = 32'd65; 
32'd1716: dataIn2 = 32'd60; 
32'd1717: dataIn2 = 32'd38; 
32'd1718: dataIn2 = 32'd77; 
32'd1719: dataIn2 = 32'd84; 
32'd1720: dataIn2 = 32'd21; 
32'd1721: dataIn2 = 32'd94; 
32'd1722: dataIn2 = 32'd63; 
32'd1723: dataIn2 = 32'd81; 
32'd1724: dataIn2 = 32'd33; 
32'd1725: dataIn2 = 32'd13; 
32'd1726: dataIn2 = 32'd46; 
32'd1727: dataIn2 = 32'd76; 
32'd1728: dataIn2 = 32'd72; 
32'd1729: dataIn2 = 32'd17; 
32'd1730: dataIn2 = 32'd79; 
32'd1731: dataIn2 = 32'd62; 
32'd1732: dataIn2 = 32'd17; 
32'd1733: dataIn2 = 32'd35; 
32'd1734: dataIn2 = 32'd79; 
32'd1735: dataIn2 = 32'd79; 
32'd1736: dataIn2 = 32'd64; 
32'd1737: dataIn2 = 32'd76; 
32'd1738: dataIn2 = 32'd27; 
32'd1739: dataIn2 = 32'd68; 
32'd1740: dataIn2 = 32'd99; 
32'd1741: dataIn2 = 32'd25; 
32'd1742: dataIn2 = 32'd43; 
32'd1743: dataIn2 = 32'd70; 
32'd1744: dataIn2 = 32'd54; 
32'd1745: dataIn2 = 32'd42; 
32'd1746: dataIn2 = 32'd78; 
32'd1747: dataIn2 = 32'd0; 
32'd1748: dataIn2 = 32'd57; 
32'd1749: dataIn2 = 32'd15; 
32'd1750: dataIn2 = 32'd94; 
32'd1751: dataIn2 = 32'd28; 
32'd1752: dataIn2 = 32'd64; 
32'd1753: dataIn2 = 32'd42; 
32'd1754: dataIn2 = 32'd29; 
32'd1755: dataIn2 = 32'd88; 
32'd1756: dataIn2 = 32'd65; 
32'd1757: dataIn2 = 32'd63; 
32'd1758: dataIn2 = 32'd81; 
32'd1759: dataIn2 = 32'd91; 
32'd1760: dataIn2 = 32'd39; 
32'd1761: dataIn2 = 32'd46; 
32'd1762: dataIn2 = 32'd55; 
32'd1763: dataIn2 = 32'd15; 
32'd1764: dataIn2 = 32'd86; 
32'd1765: dataIn2 = 32'd38; 
32'd1766: dataIn2 = 32'd2; 
32'd1767: dataIn2 = 32'd21; 
32'd1768: dataIn2 = 32'd47; 
32'd1769: dataIn2 = 32'd82; 
32'd1770: dataIn2 = 32'd60; 
32'd1771: dataIn2 = 32'd54; 
32'd1772: dataIn2 = 32'd40; 
32'd1773: dataIn2 = 32'd13; 
32'd1774: dataIn2 = 32'd12; 
32'd1775: dataIn2 = 32'd76; 
32'd1776: dataIn2 = 32'd57; 
32'd1777: dataIn2 = 32'd13; 
32'd1778: dataIn2 = 32'd14; 
32'd1779: dataIn2 = 32'd10; 
32'd1780: dataIn2 = 32'd17; 
32'd1781: dataIn2 = 32'd69; 
32'd1782: dataIn2 = 32'd100; 
32'd1783: dataIn2 = 32'd35; 
32'd1784: dataIn2 = 32'd79; 
32'd1785: dataIn2 = 32'd87; 
32'd1786: dataIn2 = 32'd99; 
32'd1787: dataIn2 = 32'd83; 
32'd1788: dataIn2 = 32'd87; 
32'd1789: dataIn2 = 32'd24; 
32'd1790: dataIn2 = 32'd15; 
32'd1791: dataIn2 = 32'd79; 
32'd1792: dataIn2 = 32'd36; 
32'd1793: dataIn2 = 32'd18; 
32'd1794: dataIn2 = 32'd1; 
32'd1795: dataIn2 = 32'd4; 
32'd1796: dataIn2 = 32'd12; 
32'd1797: dataIn2 = 32'd34; 
32'd1798: dataIn2 = 32'd24; 
32'd1799: dataIn2 = 32'd83; 
32'd1800: dataIn2 = 32'd50; 
32'd1801: dataIn2 = 32'd4; 
32'd1802: dataIn2 = 32'd3; 
32'd1803: dataIn2 = 32'd49; 
32'd1804: dataIn2 = 32'd36; 
32'd1805: dataIn2 = 32'd24; 
32'd1806: dataIn2 = 32'd96; 
32'd1807: dataIn2 = 32'd70; 
32'd1808: dataIn2 = 32'd80; 
32'd1809: dataIn2 = 32'd63; 
32'd1810: dataIn2 = 32'd89; 
32'd1811: dataIn2 = 32'd10; 
32'd1812: dataIn2 = 32'd15; 
32'd1813: dataIn2 = 32'd21; 
32'd1814: dataIn2 = 32'd38; 
32'd1815: dataIn2 = 32'd54; 
32'd1816: dataIn2 = 32'd91; 
32'd1817: dataIn2 = 32'd94; 
32'd1818: dataIn2 = 32'd97; 
32'd1819: dataIn2 = 32'd17; 
32'd1820: dataIn2 = 32'd82; 
32'd1821: dataIn2 = 32'd63; 
32'd1822: dataIn2 = 32'd100; 
32'd1823: dataIn2 = 32'd73; 
32'd1824: dataIn2 = 32'd73; 
32'd1825: dataIn2 = 32'd3; 
32'd1826: dataIn2 = 32'd53; 
32'd1827: dataIn2 = 32'd25; 
32'd1828: dataIn2 = 32'd75; 
32'd1829: dataIn2 = 32'd65; 
32'd1830: dataIn2 = 32'd71; 
32'd1831: dataIn2 = 32'd82; 
32'd1832: dataIn2 = 32'd64; 
32'd1833: dataIn2 = 32'd74; 
32'd1834: dataIn2 = 32'd10; 
32'd1835: dataIn2 = 32'd59; 
32'd1836: dataIn2 = 32'd82; 
32'd1837: dataIn2 = 32'd51; 
32'd1838: dataIn2 = 32'd59; 
32'd1839: dataIn2 = 32'd62; 
32'd1840: dataIn2 = 32'd49; 
32'd1841: dataIn2 = 32'd34; 
32'd1842: dataIn2 = 32'd39; 
32'd1843: dataIn2 = 32'd80; 
32'd1844: dataIn2 = 32'd91; 
32'd1845: dataIn2 = 32'd23; 
32'd1846: dataIn2 = 32'd40; 
32'd1847: dataIn2 = 32'd20; 
32'd1848: dataIn2 = 32'd47; 
32'd1849: dataIn2 = 32'd98; 
32'd1850: dataIn2 = 32'd86; 
32'd1851: dataIn2 = 32'd69; 
32'd1852: dataIn2 = 32'd94; 
32'd1853: dataIn2 = 32'd28; 
32'd1854: dataIn2 = 32'd19; 
32'd1855: dataIn2 = 32'd80; 
32'd1856: dataIn2 = 32'd65; 
32'd1857: dataIn2 = 32'd96; 
32'd1858: dataIn2 = 32'd28; 
32'd1859: dataIn2 = 32'd16; 
32'd1860: dataIn2 = 32'd92; 
32'd1861: dataIn2 = 32'd42; 
32'd1862: dataIn2 = 32'd27; 
32'd1863: dataIn2 = 32'd72; 
32'd1864: dataIn2 = 32'd45; 
32'd1865: dataIn2 = 32'd51; 
32'd1866: dataIn2 = 32'd2; 
32'd1867: dataIn2 = 32'd58; 
32'd1868: dataIn2 = 32'd61; 
32'd1869: dataIn2 = 32'd6; 
32'd1870: dataIn2 = 32'd40; 
32'd1871: dataIn2 = 32'd79; 
32'd1872: dataIn2 = 32'd67; 
32'd1873: dataIn2 = 32'd31; 
32'd1874: dataIn2 = 32'd19; 
32'd1875: dataIn2 = 32'd67; 
32'd1876: dataIn2 = 32'd0; 
32'd1877: dataIn2 = 32'd90; 
32'd1878: dataIn2 = 32'd29; 
32'd1879: dataIn2 = 32'd26; 
32'd1880: dataIn2 = 32'd94; 
32'd1881: dataIn2 = 32'd97; 
32'd1882: dataIn2 = 32'd40; 
32'd1883: dataIn2 = 32'd55; 
32'd1884: dataIn2 = 32'd14; 
32'd1885: dataIn2 = 32'd83; 
32'd1886: dataIn2 = 32'd5; 
32'd1887: dataIn2 = 32'd4; 
32'd1888: dataIn2 = 32'd59; 
32'd1889: dataIn2 = 32'd95; 
32'd1890: dataIn2 = 32'd32; 
32'd1891: dataIn2 = 32'd27; 
32'd1892: dataIn2 = 32'd79; 
32'd1893: dataIn2 = 32'd70; 
32'd1894: dataIn2 = 32'd57; 
32'd1895: dataIn2 = 32'd19; 
32'd1896: dataIn2 = 32'd70; 
32'd1897: dataIn2 = 32'd79; 
32'd1898: dataIn2 = 32'd40; 
32'd1899: dataIn2 = 32'd70; 
32'd1900: dataIn2 = 32'd2; 
32'd1901: dataIn2 = 32'd13; 
32'd1902: dataIn2 = 32'd6; 
32'd1903: dataIn2 = 32'd90; 
32'd1904: dataIn2 = 32'd72; 
32'd1905: dataIn2 = 32'd15; 
32'd1906: dataIn2 = 32'd46; 
32'd1907: dataIn2 = 32'd94; 
32'd1908: dataIn2 = 32'd90; 
32'd1909: dataIn2 = 32'd8; 
32'd1910: dataIn2 = 32'd78; 
32'd1911: dataIn2 = 32'd80; 
32'd1912: dataIn2 = 32'd45; 
32'd1913: dataIn2 = 32'd76; 
32'd1914: dataIn2 = 32'd23; 
32'd1915: dataIn2 = 32'd91; 
32'd1916: dataIn2 = 32'd2; 
32'd1917: dataIn2 = 32'd80; 
32'd1918: dataIn2 = 32'd21; 
32'd1919: dataIn2 = 32'd36; 
32'd1920: dataIn2 = 32'd17; 
32'd1921: dataIn2 = 32'd14; 
32'd1922: dataIn2 = 32'd78; 
32'd1923: dataIn2 = 32'd41; 
32'd1924: dataIn2 = 32'd68; 
32'd1925: dataIn2 = 32'd54; 
32'd1926: dataIn2 = 32'd35; 
32'd1927: dataIn2 = 32'd59; 
32'd1928: dataIn2 = 32'd71; 
32'd1929: dataIn2 = 32'd74; 
32'd1930: dataIn2 = 32'd22; 
32'd1931: dataIn2 = 32'd80; 
32'd1932: dataIn2 = 32'd47; 
32'd1933: dataIn2 = 32'd76; 
32'd1934: dataIn2 = 32'd5; 
32'd1935: dataIn2 = 32'd2; 
32'd1936: dataIn2 = 32'd71; 
32'd1937: dataIn2 = 32'd1; 
32'd1938: dataIn2 = 32'd13; 
32'd1939: dataIn2 = 32'd55; 
32'd1940: dataIn2 = 32'd81; 
32'd1941: dataIn2 = 32'd27; 
32'd1942: dataIn2 = 32'd66; 
32'd1943: dataIn2 = 32'd63; 
32'd1944: dataIn2 = 32'd47; 
32'd1945: dataIn2 = 32'd17; 
32'd1946: dataIn2 = 32'd6; 
32'd1947: dataIn2 = 32'd91; 
32'd1948: dataIn2 = 32'd24; 
32'd1949: dataIn2 = 32'd48; 
32'd1950: dataIn2 = 32'd0; 
32'd1951: dataIn2 = 32'd96; 
32'd1952: dataIn2 = 32'd48; 
32'd1953: dataIn2 = 32'd25; 
32'd1954: dataIn2 = 32'd2; 
32'd1955: dataIn2 = 32'd77; 
32'd1956: dataIn2 = 32'd43; 
32'd1957: dataIn2 = 32'd29; 
32'd1958: dataIn2 = 32'd10; 
32'd1959: dataIn2 = 32'd96; 
32'd1960: dataIn2 = 32'd35; 
32'd1961: dataIn2 = 32'd90; 
32'd1962: dataIn2 = 32'd34; 
32'd1963: dataIn2 = 32'd2; 
32'd1964: dataIn2 = 32'd47; 
32'd1965: dataIn2 = 32'd22; 
32'd1966: dataIn2 = 32'd99; 
32'd1967: dataIn2 = 32'd86; 
32'd1968: dataIn2 = 32'd85; 
32'd1969: dataIn2 = 32'd17; 
32'd1970: dataIn2 = 32'd34; 
32'd1971: dataIn2 = 32'd17; 
32'd1972: dataIn2 = 32'd69; 
32'd1973: dataIn2 = 32'd13; 
32'd1974: dataIn2 = 32'd11; 
32'd1975: dataIn2 = 32'd34; 
32'd1976: dataIn2 = 32'd52; 
32'd1977: dataIn2 = 32'd39; 
32'd1978: dataIn2 = 32'd38; 
32'd1979: dataIn2 = 32'd6; 
32'd1980: dataIn2 = 32'd77; 
32'd1981: dataIn2 = 32'd80; 
32'd1982: dataIn2 = 32'd26; 
32'd1983: dataIn2 = 32'd7; 
32'd1984: dataIn2 = 32'd44; 
32'd1985: dataIn2 = 32'd87; 
32'd1986: dataIn2 = 32'd97; 
32'd1987: dataIn2 = 32'd79; 
32'd1988: dataIn2 = 32'd77; 
32'd1989: dataIn2 = 32'd45; 
32'd1990: dataIn2 = 32'd16; 
32'd1991: dataIn2 = 32'd8; 
32'd1992: dataIn2 = 32'd24; 
32'd1993: dataIn2 = 32'd11; 
32'd1994: dataIn2 = 32'd27; 
32'd1995: dataIn2 = 32'd88; 
32'd1996: dataIn2 = 32'd90; 
32'd1997: dataIn2 = 32'd8; 
32'd1998: dataIn2 = 32'd36; 
32'd1999: dataIn2 = 32'd9; 
32'd2000: dataIn2 = 32'd26; 
32'd2001: dataIn2 = 32'd74; 
32'd2002: dataIn2 = 32'd68; 
32'd2003: dataIn2 = 32'd89; 
32'd2004: dataIn2 = 32'd35; 
32'd2005: dataIn2 = 32'd70; 
32'd2006: dataIn2 = 32'd97; 
32'd2007: dataIn2 = 32'd44; 
32'd2008: dataIn2 = 32'd29; 
32'd2009: dataIn2 = 32'd23; 
32'd2010: dataIn2 = 32'd42; 
32'd2011: dataIn2 = 32'd18; 
32'd2012: dataIn2 = 32'd92; 
32'd2013: dataIn2 = 32'd6; 
32'd2014: dataIn2 = 32'd67; 
32'd2015: dataIn2 = 32'd6; 
32'd2016: dataIn2 = 32'd87; 
32'd2017: dataIn2 = 32'd49; 
32'd2018: dataIn2 = 32'd54; 
32'd2019: dataIn2 = 32'd79; 
32'd2020: dataIn2 = 32'd13; 
32'd2021: dataIn2 = 32'd22; 
32'd2022: dataIn2 = 32'd2; 
32'd2023: dataIn2 = 32'd84; 
32'd2024: dataIn2 = 32'd13; 
32'd2025: dataIn2 = 32'd2; 
32'd2026: dataIn2 = 32'd63; 
32'd2027: dataIn2 = 32'd52; 
32'd2028: dataIn2 = 32'd34; 
32'd2029: dataIn2 = 32'd61; 
32'd2030: dataIn2 = 32'd82; 
32'd2031: dataIn2 = 32'd76; 
32'd2032: dataIn2 = 32'd45; 
32'd2033: dataIn2 = 32'd39; 
32'd2034: dataIn2 = 32'd16; 
32'd2035: dataIn2 = 32'd46; 
32'd2036: dataIn2 = 32'd80; 
32'd2037: dataIn2 = 32'd72; 
32'd2038: dataIn2 = 32'd63; 
32'd2039: dataIn2 = 32'd48; 
32'd2040: dataIn2 = 32'd27; 
32'd2041: dataIn2 = 32'd100; 
32'd2042: dataIn2 = 32'd75; 
32'd2043: dataIn2 = 32'd67; 
32'd2044: dataIn2 = 32'd5; 
32'd2045: dataIn2 = 32'd42; 
32'd2046: dataIn2 = 32'd95; 
32'd2047: dataIn2 = 32'd86; 
32'd2048: dataIn2 = 32'd49; 
32'd2049: dataIn2 = 32'd61; 
32'd2050: dataIn2 = 32'd59; 
32'd2051: dataIn2 = 32'd62; 
32'd2052: dataIn2 = 32'd71; 
32'd2053: dataIn2 = 32'd58; 
32'd2054: dataIn2 = 32'd53; 
32'd2055: dataIn2 = 32'd17; 
32'd2056: dataIn2 = 32'd99; 
32'd2057: dataIn2 = 32'd60; 
32'd2058: dataIn2 = 32'd27; 
32'd2059: dataIn2 = 32'd98; 
32'd2060: dataIn2 = 32'd6; 
32'd2061: dataIn2 = 32'd58; 
32'd2062: dataIn2 = 32'd48; 
32'd2063: dataIn2 = 32'd76; 
32'd2064: dataIn2 = 32'd42; 
32'd2065: dataIn2 = 32'd72; 
32'd2066: dataIn2 = 32'd10; 
32'd2067: dataIn2 = 32'd9; 
32'd2068: dataIn2 = 32'd78; 
32'd2069: dataIn2 = 32'd23; 
32'd2070: dataIn2 = 32'd65; 
32'd2071: dataIn2 = 32'd70; 
32'd2072: dataIn2 = 32'd89; 
32'd2073: dataIn2 = 32'd54; 
32'd2074: dataIn2 = 32'd35; 
32'd2075: dataIn2 = 32'd5; 
32'd2076: dataIn2 = 32'd67; 
32'd2077: dataIn2 = 32'd19; 
32'd2078: dataIn2 = 32'd66; 
32'd2079: dataIn2 = 32'd1; 
32'd2080: dataIn2 = 32'd87; 
32'd2081: dataIn2 = 32'd95; 
32'd2082: dataIn2 = 32'd61; 
32'd2083: dataIn2 = 32'd76; 
32'd2084: dataIn2 = 32'd49; 
32'd2085: dataIn2 = 32'd27; 
32'd2086: dataIn2 = 32'd14; 
32'd2087: dataIn2 = 32'd66; 
32'd2088: dataIn2 = 32'd12; 
32'd2089: dataIn2 = 32'd16; 
32'd2090: dataIn2 = 32'd80; 
32'd2091: dataIn2 = 32'd93; 
32'd2092: dataIn2 = 32'd62; 
32'd2093: dataIn2 = 32'd88; 
32'd2094: dataIn2 = 32'd41; 
32'd2095: dataIn2 = 32'd92; 
32'd2096: dataIn2 = 32'd38; 
32'd2097: dataIn2 = 32'd43; 
32'd2098: dataIn2 = 32'd74; 
32'd2099: dataIn2 = 32'd24; 
32'd2100: dataIn2 = 32'd75; 
32'd2101: dataIn2 = 32'd49; 
32'd2102: dataIn2 = 32'd20; 
32'd2103: dataIn2 = 32'd86; 
32'd2104: dataIn2 = 32'd13; 
32'd2105: dataIn2 = 32'd60; 
32'd2106: dataIn2 = 32'd28; 
32'd2107: dataIn2 = 32'd100; 
32'd2108: dataIn2 = 32'd21; 
32'd2109: dataIn2 = 32'd68; 
32'd2110: dataIn2 = 32'd57; 
32'd2111: dataIn2 = 32'd22; 
32'd2112: dataIn2 = 32'd36; 
32'd2113: dataIn2 = 32'd30; 
32'd2114: dataIn2 = 32'd11; 
32'd2115: dataIn2 = 32'd97; 
32'd2116: dataIn2 = 32'd84; 
32'd2117: dataIn2 = 32'd48; 
32'd2118: dataIn2 = 32'd30; 
32'd2119: dataIn2 = 32'd2; 
32'd2120: dataIn2 = 32'd31; 
32'd2121: dataIn2 = 32'd35; 
32'd2122: dataIn2 = 32'd61; 
32'd2123: dataIn2 = 32'd64; 
32'd2124: dataIn2 = 32'd77; 
32'd2125: dataIn2 = 32'd30; 
32'd2126: dataIn2 = 32'd16; 
32'd2127: dataIn2 = 32'd10; 
32'd2128: dataIn2 = 32'd82; 
32'd2129: dataIn2 = 32'd15; 
32'd2130: dataIn2 = 32'd100; 
32'd2131: dataIn2 = 32'd43; 
32'd2132: dataIn2 = 32'd69; 
32'd2133: dataIn2 = 32'd79; 
32'd2134: dataIn2 = 32'd33; 
32'd2135: dataIn2 = 32'd94; 
32'd2136: dataIn2 = 32'd65; 
32'd2137: dataIn2 = 32'd83; 
32'd2138: dataIn2 = 32'd97; 
32'd2139: dataIn2 = 32'd63; 
32'd2140: dataIn2 = 32'd15; 
32'd2141: dataIn2 = 32'd49; 
32'd2142: dataIn2 = 32'd35; 
32'd2143: dataIn2 = 32'd0; 
32'd2144: dataIn2 = 32'd4; 
32'd2145: dataIn2 = 32'd38; 
32'd2146: dataIn2 = 32'd46; 
32'd2147: dataIn2 = 32'd69; 
32'd2148: dataIn2 = 32'd92; 
32'd2149: dataIn2 = 32'd35; 
32'd2150: dataIn2 = 32'd4; 
32'd2151: dataIn2 = 32'd42; 
32'd2152: dataIn2 = 32'd58; 
32'd2153: dataIn2 = 32'd62; 
32'd2154: dataIn2 = 32'd17; 
32'd2155: dataIn2 = 32'd51; 
32'd2156: dataIn2 = 32'd50; 
32'd2157: dataIn2 = 32'd18; 
32'd2158: dataIn2 = 32'd68; 
32'd2159: dataIn2 = 32'd93; 
32'd2160: dataIn2 = 32'd42; 
32'd2161: dataIn2 = 32'd12; 
32'd2162: dataIn2 = 32'd56; 
32'd2163: dataIn2 = 32'd23; 
32'd2164: dataIn2 = 32'd18; 
32'd2165: dataIn2 = 32'd19; 
32'd2166: dataIn2 = 32'd45; 
32'd2167: dataIn2 = 32'd1; 
32'd2168: dataIn2 = 32'd72; 
32'd2169: dataIn2 = 32'd95; 
32'd2170: dataIn2 = 32'd30; 
32'd2171: dataIn2 = 32'd32; 
32'd2172: dataIn2 = 32'd38; 
32'd2173: dataIn2 = 32'd49; 
32'd2174: dataIn2 = 32'd51; 
32'd2175: dataIn2 = 32'd23; 
32'd2176: dataIn2 = 32'd96; 
32'd2177: dataIn2 = 32'd63; 
32'd2178: dataIn2 = 32'd52; 
32'd2179: dataIn2 = 32'd32; 
32'd2180: dataIn2 = 32'd53; 
32'd2181: dataIn2 = 32'd38; 
32'd2182: dataIn2 = 32'd11; 
32'd2183: dataIn2 = 32'd90; 
32'd2184: dataIn2 = 32'd56; 
32'd2185: dataIn2 = 32'd69; 
32'd2186: dataIn2 = 32'd75; 
32'd2187: dataIn2 = 32'd48; 
32'd2188: dataIn2 = 32'd98; 
32'd2189: dataIn2 = 32'd45; 
32'd2190: dataIn2 = 32'd98; 
32'd2191: dataIn2 = 32'd28; 
32'd2192: dataIn2 = 32'd7; 
32'd2193: dataIn2 = 32'd25; 
32'd2194: dataIn2 = 32'd74; 
32'd2195: dataIn2 = 32'd97; 
32'd2196: dataIn2 = 32'd7; 
32'd2197: dataIn2 = 32'd37; 
32'd2198: dataIn2 = 32'd39; 
32'd2199: dataIn2 = 32'd38; 
32'd2200: dataIn2 = 32'd74; 
32'd2201: dataIn2 = 32'd4; 
32'd2202: dataIn2 = 32'd6; 
32'd2203: dataIn2 = 32'd54; 
32'd2204: dataIn2 = 32'd42; 
32'd2205: dataIn2 = 32'd88; 
32'd2206: dataIn2 = 32'd68; 
32'd2207: dataIn2 = 32'd52; 
32'd2208: dataIn2 = 32'd17; 
32'd2209: dataIn2 = 32'd69; 
32'd2210: dataIn2 = 32'd71; 
32'd2211: dataIn2 = 32'd7; 
32'd2212: dataIn2 = 32'd100; 
32'd2213: dataIn2 = 32'd32; 
32'd2214: dataIn2 = 32'd49; 
32'd2215: dataIn2 = 32'd57; 
32'd2216: dataIn2 = 32'd24; 
32'd2217: dataIn2 = 32'd53; 
32'd2218: dataIn2 = 32'd25; 
32'd2219: dataIn2 = 32'd6; 
32'd2220: dataIn2 = 32'd63; 
32'd2221: dataIn2 = 32'd88; 
32'd2222: dataIn2 = 32'd94; 
32'd2223: dataIn2 = 32'd90; 
32'd2224: dataIn2 = 32'd0; 
32'd2225: dataIn2 = 32'd40; 
32'd2226: dataIn2 = 32'd66; 
32'd2227: dataIn2 = 32'd34; 
32'd2228: dataIn2 = 32'd27; 
32'd2229: dataIn2 = 32'd41; 
32'd2230: dataIn2 = 32'd56; 
32'd2231: dataIn2 = 32'd7; 
32'd2232: dataIn2 = 32'd77; 
32'd2233: dataIn2 = 32'd47; 
32'd2234: dataIn2 = 32'd23; 
32'd2235: dataIn2 = 32'd31; 
32'd2236: dataIn2 = 32'd50; 
32'd2237: dataIn2 = 32'd17; 
32'd2238: dataIn2 = 32'd1; 
32'd2239: dataIn2 = 32'd34; 
32'd2240: dataIn2 = 32'd86; 
32'd2241: dataIn2 = 32'd34; 
32'd2242: dataIn2 = 32'd64; 
32'd2243: dataIn2 = 32'd25; 
32'd2244: dataIn2 = 32'd30; 
32'd2245: dataIn2 = 32'd57; 
32'd2246: dataIn2 = 32'd32; 
32'd2247: dataIn2 = 32'd12; 
32'd2248: dataIn2 = 32'd83; 
32'd2249: dataIn2 = 32'd24; 
32'd2250: dataIn2 = 32'd78; 
32'd2251: dataIn2 = 32'd22; 
32'd2252: dataIn2 = 32'd81; 
32'd2253: dataIn2 = 32'd73; 
32'd2254: dataIn2 = 32'd35; 
32'd2255: dataIn2 = 32'd65; 
32'd2256: dataIn2 = 32'd99; 
32'd2257: dataIn2 = 32'd20; 
32'd2258: dataIn2 = 32'd15; 
32'd2259: dataIn2 = 32'd47; 
32'd2260: dataIn2 = 32'd29; 
32'd2261: dataIn2 = 32'd16; 
32'd2262: dataIn2 = 32'd12; 
32'd2263: dataIn2 = 32'd69; 
32'd2264: dataIn2 = 32'd90; 
32'd2265: dataIn2 = 32'd92; 
32'd2266: dataIn2 = 32'd65; 
32'd2267: dataIn2 = 32'd26; 
32'd2268: dataIn2 = 32'd3; 
32'd2269: dataIn2 = 32'd4; 
32'd2270: dataIn2 = 32'd79; 
32'd2271: dataIn2 = 32'd98; 
32'd2272: dataIn2 = 32'd44; 
32'd2273: dataIn2 = 32'd34; 
32'd2274: dataIn2 = 32'd95; 
32'd2275: dataIn2 = 32'd15; 
32'd2276: dataIn2 = 32'd48; 
32'd2277: dataIn2 = 32'd36; 
32'd2278: dataIn2 = 32'd4; 
32'd2279: dataIn2 = 32'd20; 
32'd2280: dataIn2 = 32'd54; 
32'd2281: dataIn2 = 32'd100; 
32'd2282: dataIn2 = 32'd98; 
32'd2283: dataIn2 = 32'd88; 
32'd2284: dataIn2 = 32'd94; 
32'd2285: dataIn2 = 32'd45; 
32'd2286: dataIn2 = 32'd28; 
32'd2287: dataIn2 = 32'd38; 
32'd2288: dataIn2 = 32'd100; 
32'd2289: dataIn2 = 32'd13; 
32'd2290: dataIn2 = 32'd42; 
32'd2291: dataIn2 = 32'd22; 
32'd2292: dataIn2 = 32'd16; 
32'd2293: dataIn2 = 32'd9; 
32'd2294: dataIn2 = 32'd6; 
32'd2295: dataIn2 = 32'd36; 
32'd2296: dataIn2 = 32'd18; 
32'd2297: dataIn2 = 32'd27; 
32'd2298: dataIn2 = 32'd75; 
32'd2299: dataIn2 = 32'd89; 
32'd2300: dataIn2 = 32'd51; 
32'd2301: dataIn2 = 32'd24; 
32'd2302: dataIn2 = 32'd30; 
32'd2303: dataIn2 = 32'd62; 
32'd2304: dataIn2 = 32'd17; 
32'd2305: dataIn2 = 32'd1; 
32'd2306: dataIn2 = 32'd45; 
32'd2307: dataIn2 = 32'd60; 
32'd2308: dataIn2 = 32'd90; 
32'd2309: dataIn2 = 32'd6; 
32'd2310: dataIn2 = 32'd82; 
32'd2311: dataIn2 = 32'd83; 
32'd2312: dataIn2 = 32'd1; 
32'd2313: dataIn2 = 32'd5; 
32'd2314: dataIn2 = 32'd33; 
32'd2315: dataIn2 = 32'd20; 
32'd2316: dataIn2 = 32'd58; 
32'd2317: dataIn2 = 32'd48; 
32'd2318: dataIn2 = 32'd31; 
32'd2319: dataIn2 = 32'd23; 
32'd2320: dataIn2 = 32'd26; 
32'd2321: dataIn2 = 32'd24; 
32'd2322: dataIn2 = 32'd88; 
32'd2323: dataIn2 = 32'd14; 
32'd2324: dataIn2 = 32'd56; 
32'd2325: dataIn2 = 32'd19; 
32'd2326: dataIn2 = 32'd28; 
32'd2327: dataIn2 = 32'd79; 
32'd2328: dataIn2 = 32'd2; 
32'd2329: dataIn2 = 32'd76; 
32'd2330: dataIn2 = 32'd3; 
32'd2331: dataIn2 = 32'd89; 
32'd2332: dataIn2 = 32'd5; 
32'd2333: dataIn2 = 32'd67; 
32'd2334: dataIn2 = 32'd40; 
32'd2335: dataIn2 = 32'd38; 
32'd2336: dataIn2 = 32'd82; 
32'd2337: dataIn2 = 32'd38; 
32'd2338: dataIn2 = 32'd13; 
32'd2339: dataIn2 = 32'd58; 
32'd2340: dataIn2 = 32'd33; 
32'd2341: dataIn2 = 32'd29; 
32'd2342: dataIn2 = 32'd21; 
32'd2343: dataIn2 = 32'd3; 
32'd2344: dataIn2 = 32'd27; 
32'd2345: dataIn2 = 32'd35; 
32'd2346: dataIn2 = 32'd90; 
32'd2347: dataIn2 = 32'd44; 
32'd2348: dataIn2 = 32'd27; 
32'd2349: dataIn2 = 32'd24; 
32'd2350: dataIn2 = 32'd1; 
32'd2351: dataIn2 = 32'd91; 
32'd2352: dataIn2 = 32'd76; 
32'd2353: dataIn2 = 32'd2; 
32'd2354: dataIn2 = 32'd36; 
32'd2355: dataIn2 = 32'd100; 
32'd2356: dataIn2 = 32'd60; 
32'd2357: dataIn2 = 32'd51; 
32'd2358: dataIn2 = 32'd86; 
32'd2359: dataIn2 = 32'd74; 
32'd2360: dataIn2 = 32'd84; 
32'd2361: dataIn2 = 32'd76; 
32'd2362: dataIn2 = 32'd41; 
32'd2363: dataIn2 = 32'd14; 
32'd2364: dataIn2 = 32'd23; 
32'd2365: dataIn2 = 32'd12; 
32'd2366: dataIn2 = 32'd82; 
32'd2367: dataIn2 = 32'd17; 
32'd2368: dataIn2 = 32'd33; 
32'd2369: dataIn2 = 32'd95; 
32'd2370: dataIn2 = 32'd66; 
32'd2371: dataIn2 = 32'd49; 
32'd2372: dataIn2 = 32'd25; 
32'd2373: dataIn2 = 32'd60; 
32'd2374: dataIn2 = 32'd6; 
32'd2375: dataIn2 = 32'd80; 
32'd2376: dataIn2 = 32'd87; 
32'd2377: dataIn2 = 32'd40; 
32'd2378: dataIn2 = 32'd21; 
32'd2379: dataIn2 = 32'd11; 
32'd2380: dataIn2 = 32'd53; 
32'd2381: dataIn2 = 32'd99; 
32'd2382: dataIn2 = 32'd78; 
32'd2383: dataIn2 = 32'd93; 
32'd2384: dataIn2 = 32'd75; 
32'd2385: dataIn2 = 32'd61; 
32'd2386: dataIn2 = 32'd69; 
32'd2387: dataIn2 = 32'd29; 
32'd2388: dataIn2 = 32'd13; 
32'd2389: dataIn2 = 32'd17; 
32'd2390: dataIn2 = 32'd100; 
32'd2391: dataIn2 = 32'd2; 
32'd2392: dataIn2 = 32'd7; 
32'd2393: dataIn2 = 32'd12; 
32'd2394: dataIn2 = 32'd99; 
32'd2395: dataIn2 = 32'd20; 
32'd2396: dataIn2 = 32'd36; 
32'd2397: dataIn2 = 32'd18; 
32'd2398: dataIn2 = 32'd20; 
32'd2399: dataIn2 = 32'd90; 
32'd2400: dataIn2 = 32'd3; 
32'd2401: dataIn2 = 32'd39; 
32'd2402: dataIn2 = 32'd54; 
32'd2403: dataIn2 = 32'd55; 
32'd2404: dataIn2 = 32'd78; 
32'd2405: dataIn2 = 32'd26; 
32'd2406: dataIn2 = 32'd97; 
32'd2407: dataIn2 = 32'd36; 
32'd2408: dataIn2 = 32'd86; 
32'd2409: dataIn2 = 32'd34; 
32'd2410: dataIn2 = 32'd7; 
32'd2411: dataIn2 = 32'd25; 
32'd2412: dataIn2 = 32'd29; 
32'd2413: dataIn2 = 32'd81; 
32'd2414: dataIn2 = 32'd20; 
32'd2415: dataIn2 = 32'd78; 
32'd2416: dataIn2 = 32'd33; 
32'd2417: dataIn2 = 32'd36; 
32'd2418: dataIn2 = 32'd62; 
32'd2419: dataIn2 = 32'd16; 
32'd2420: dataIn2 = 32'd3; 
32'd2421: dataIn2 = 32'd91; 
32'd2422: dataIn2 = 32'd53; 
32'd2423: dataIn2 = 32'd22; 
32'd2424: dataIn2 = 32'd84; 
32'd2425: dataIn2 = 32'd40; 
32'd2426: dataIn2 = 32'd95; 
32'd2427: dataIn2 = 32'd11; 
32'd2428: dataIn2 = 32'd92; 
32'd2429: dataIn2 = 32'd62; 
32'd2430: dataIn2 = 32'd73; 
32'd2431: dataIn2 = 32'd2; 
32'd2432: dataIn2 = 32'd77; 
32'd2433: dataIn2 = 32'd95; 
32'd2434: dataIn2 = 32'd40; 
32'd2435: dataIn2 = 32'd76; 
32'd2436: dataIn2 = 32'd100; 
32'd2437: dataIn2 = 32'd49; 
32'd2438: dataIn2 = 32'd83; 
32'd2439: dataIn2 = 32'd48; 
32'd2440: dataIn2 = 32'd91; 
32'd2441: dataIn2 = 32'd26; 
32'd2442: dataIn2 = 32'd98; 
32'd2443: dataIn2 = 32'd77; 
32'd2444: dataIn2 = 32'd19; 
32'd2445: dataIn2 = 32'd86; 
32'd2446: dataIn2 = 32'd95; 
32'd2447: dataIn2 = 32'd47; 
32'd2448: dataIn2 = 32'd24; 
32'd2449: dataIn2 = 32'd16; 
32'd2450: dataIn2 = 32'd1; 
32'd2451: dataIn2 = 32'd25; 
32'd2452: dataIn2 = 32'd10; 
32'd2453: dataIn2 = 32'd81; 
32'd2454: dataIn2 = 32'd8; 
32'd2455: dataIn2 = 32'd16; 
32'd2456: dataIn2 = 32'd10; 
32'd2457: dataIn2 = 32'd14; 
32'd2458: dataIn2 = 32'd0; 
32'd2459: dataIn2 = 32'd32; 
32'd2460: dataIn2 = 32'd80; 
32'd2461: dataIn2 = 32'd60; 
32'd2462: dataIn2 = 32'd31; 
32'd2463: dataIn2 = 32'd85; 
32'd2464: dataIn2 = 32'd43; 
32'd2465: dataIn2 = 32'd90; 
32'd2466: dataIn2 = 32'd74; 
32'd2467: dataIn2 = 32'd58; 
32'd2468: dataIn2 = 32'd5; 
32'd2469: dataIn2 = 32'd41; 
32'd2470: dataIn2 = 32'd30; 
32'd2471: dataIn2 = 32'd21; 
32'd2472: dataIn2 = 32'd61; 
32'd2473: dataIn2 = 32'd20; 
32'd2474: dataIn2 = 32'd94; 
32'd2475: dataIn2 = 32'd59; 
32'd2476: dataIn2 = 32'd94; 
32'd2477: dataIn2 = 32'd25; 
32'd2478: dataIn2 = 32'd28; 
32'd2479: dataIn2 = 32'd50; 
32'd2480: dataIn2 = 32'd63; 
32'd2481: dataIn2 = 32'd86; 
32'd2482: dataIn2 = 32'd63; 
32'd2483: dataIn2 = 32'd70; 
32'd2484: dataIn2 = 32'd93; 
32'd2485: dataIn2 = 32'd48; 
32'd2486: dataIn2 = 32'd46; 
32'd2487: dataIn2 = 32'd4; 
32'd2488: dataIn2 = 32'd31; 
32'd2489: dataIn2 = 32'd29; 
32'd2490: dataIn2 = 32'd50; 
32'd2491: dataIn2 = 32'd68; 
32'd2492: dataIn2 = 32'd54; 
32'd2493: dataIn2 = 32'd88; 
32'd2494: dataIn2 = 32'd92; 
32'd2495: dataIn2 = 32'd65; 
32'd2496: dataIn2 = 32'd71; 
32'd2497: dataIn2 = 32'd60; 
32'd2498: dataIn2 = 32'd15; 
32'd2499: dataIn2 = 32'd81; 
32'd2500: dataIn2 = 32'd59; 
32'd2501: dataIn2 = 32'd8; 
32'd2502: dataIn2 = 32'd92; 
32'd2503: dataIn2 = 32'd55; 
32'd2504: dataIn2 = 32'd88; 
32'd2505: dataIn2 = 32'd40; 
32'd2506: dataIn2 = 32'd47; 
32'd2507: dataIn2 = 32'd50; 
32'd2508: dataIn2 = 32'd95; 
32'd2509: dataIn2 = 32'd12; 
32'd2510: dataIn2 = 32'd100; 
32'd2511: dataIn2 = 32'd19; 
32'd2512: dataIn2 = 32'd32; 
32'd2513: dataIn2 = 32'd9; 
32'd2514: dataIn2 = 32'd17; 
32'd2515: dataIn2 = 32'd89; 
32'd2516: dataIn2 = 32'd93; 
32'd2517: dataIn2 = 32'd95; 
32'd2518: dataIn2 = 32'd75; 
32'd2519: dataIn2 = 32'd75; 
32'd2520: dataIn2 = 32'd93; 
32'd2521: dataIn2 = 32'd84; 
32'd2522: dataIn2 = 32'd41; 
32'd2523: dataIn2 = 32'd95; 
32'd2524: dataIn2 = 32'd40; 
32'd2525: dataIn2 = 32'd30; 
32'd2526: dataIn2 = 32'd89; 
32'd2527: dataIn2 = 32'd28; 
32'd2528: dataIn2 = 32'd87; 
32'd2529: dataIn2 = 32'd89; 
32'd2530: dataIn2 = 32'd47; 
32'd2531: dataIn2 = 32'd89; 
32'd2532: dataIn2 = 32'd85; 
32'd2533: dataIn2 = 32'd21; 
32'd2534: dataIn2 = 32'd86; 
32'd2535: dataIn2 = 32'd75; 
32'd2536: dataIn2 = 32'd26; 
32'd2537: dataIn2 = 32'd32; 
32'd2538: dataIn2 = 32'd91; 
32'd2539: dataIn2 = 32'd56; 
32'd2540: dataIn2 = 32'd78; 
32'd2541: dataIn2 = 32'd70; 
32'd2542: dataIn2 = 32'd2; 
32'd2543: dataIn2 = 32'd51; 
32'd2544: dataIn2 = 32'd63; 
32'd2545: dataIn2 = 32'd70; 
32'd2546: dataIn2 = 32'd15; 
32'd2547: dataIn2 = 32'd76; 
32'd2548: dataIn2 = 32'd41; 
32'd2549: dataIn2 = 32'd90; 
32'd2550: dataIn2 = 32'd20; 
32'd2551: dataIn2 = 32'd84; 
32'd2552: dataIn2 = 32'd98; 
32'd2553: dataIn2 = 32'd93; 
32'd2554: dataIn2 = 32'd3; 
32'd2555: dataIn2 = 32'd56; 
32'd2556: dataIn2 = 32'd70; 
32'd2557: dataIn2 = 32'd23; 
32'd2558: dataIn2 = 32'd20; 
32'd2559: dataIn2 = 32'd51; 
32'd2560: dataIn2 = 32'd78; 
32'd2561: dataIn2 = 32'd62; 
32'd2562: dataIn2 = 32'd31; 
32'd2563: dataIn2 = 32'd21; 
32'd2564: dataIn2 = 32'd61; 
32'd2565: dataIn2 = 32'd5; 
32'd2566: dataIn2 = 32'd57; 
32'd2567: dataIn2 = 32'd90; 
32'd2568: dataIn2 = 32'd5; 
32'd2569: dataIn2 = 32'd88; 
32'd2570: dataIn2 = 32'd78; 
32'd2571: dataIn2 = 32'd96; 
32'd2572: dataIn2 = 32'd42; 
32'd2573: dataIn2 = 32'd41; 
32'd2574: dataIn2 = 32'd73; 
32'd2575: dataIn2 = 32'd77; 
32'd2576: dataIn2 = 32'd42; 
32'd2577: dataIn2 = 32'd93; 
32'd2578: dataIn2 = 32'd41; 
32'd2579: dataIn2 = 32'd17; 
32'd2580: dataIn2 = 32'd55; 
32'd2581: dataIn2 = 32'd28; 
32'd2582: dataIn2 = 32'd33; 
32'd2583: dataIn2 = 32'd78; 
32'd2584: dataIn2 = 32'd24; 
32'd2585: dataIn2 = 32'd98; 
32'd2586: dataIn2 = 32'd15; 
32'd2587: dataIn2 = 32'd8; 
32'd2588: dataIn2 = 32'd65; 
32'd2589: dataIn2 = 32'd56; 
32'd2590: dataIn2 = 32'd58; 
32'd2591: dataIn2 = 32'd36; 
32'd2592: dataIn2 = 32'd15; 
32'd2593: dataIn2 = 32'd97; 
32'd2594: dataIn2 = 32'd56; 
32'd2595: dataIn2 = 32'd43; 
32'd2596: dataIn2 = 32'd5; 
32'd2597: dataIn2 = 32'd1; 
32'd2598: dataIn2 = 32'd46; 
32'd2599: dataIn2 = 32'd32; 
32'd2600: dataIn2 = 32'd52; 
32'd2601: dataIn2 = 32'd2; 
32'd2602: dataIn2 = 32'd89; 
32'd2603: dataIn2 = 32'd62; 
32'd2604: dataIn2 = 32'd75; 
32'd2605: dataIn2 = 32'd44; 
32'd2606: dataIn2 = 32'd56; 
32'd2607: dataIn2 = 32'd98; 
32'd2608: dataIn2 = 32'd71; 
32'd2609: dataIn2 = 32'd51; 
32'd2610: dataIn2 = 32'd76; 
32'd2611: dataIn2 = 32'd41; 
32'd2612: dataIn2 = 32'd17; 
32'd2613: dataIn2 = 32'd26; 
32'd2614: dataIn2 = 32'd5; 
32'd2615: dataIn2 = 32'd73; 
32'd2616: dataIn2 = 32'd14; 
32'd2617: dataIn2 = 32'd23; 
32'd2618: dataIn2 = 32'd56; 
32'd2619: dataIn2 = 32'd31; 
32'd2620: dataIn2 = 32'd40; 
32'd2621: dataIn2 = 32'd60; 
32'd2622: dataIn2 = 32'd48; 
32'd2623: dataIn2 = 32'd63; 
32'd2624: dataIn2 = 32'd31; 
32'd2625: dataIn2 = 32'd25; 
32'd2626: dataIn2 = 32'd31; 
32'd2627: dataIn2 = 32'd34; 
32'd2628: dataIn2 = 32'd69; 
32'd2629: dataIn2 = 32'd62; 
32'd2630: dataIn2 = 32'd39; 
32'd2631: dataIn2 = 32'd68; 
32'd2632: dataIn2 = 32'd73; 
32'd2633: dataIn2 = 32'd32; 
32'd2634: dataIn2 = 32'd100; 
32'd2635: dataIn2 = 32'd46; 
32'd2636: dataIn2 = 32'd29; 
32'd2637: dataIn2 = 32'd33; 
32'd2638: dataIn2 = 32'd55; 
32'd2639: dataIn2 = 32'd46; 
32'd2640: dataIn2 = 32'd91; 
32'd2641: dataIn2 = 32'd15; 
32'd2642: dataIn2 = 32'd53; 
32'd2643: dataIn2 = 32'd36; 
32'd2644: dataIn2 = 32'd22; 
32'd2645: dataIn2 = 32'd31; 
32'd2646: dataIn2 = 32'd86; 
32'd2647: dataIn2 = 32'd22; 
32'd2648: dataIn2 = 32'd78; 
32'd2649: dataIn2 = 32'd41; 
32'd2650: dataIn2 = 32'd22; 
32'd2651: dataIn2 = 32'd99; 
32'd2652: dataIn2 = 32'd93; 
32'd2653: dataIn2 = 32'd41; 
32'd2654: dataIn2 = 32'd33; 
32'd2655: dataIn2 = 32'd65; 
32'd2656: dataIn2 = 32'd45; 
32'd2657: dataIn2 = 32'd35; 
32'd2658: dataIn2 = 32'd18; 
32'd2659: dataIn2 = 32'd71; 
32'd2660: dataIn2 = 32'd25; 
32'd2661: dataIn2 = 32'd40; 
32'd2662: dataIn2 = 32'd41; 
32'd2663: dataIn2 = 32'd63; 
32'd2664: dataIn2 = 32'd13; 
32'd2665: dataIn2 = 32'd50; 
32'd2666: dataIn2 = 32'd3; 
32'd2667: dataIn2 = 32'd58; 
32'd2668: dataIn2 = 32'd76; 
32'd2669: dataIn2 = 32'd20; 
32'd2670: dataIn2 = 32'd58; 
32'd2671: dataIn2 = 32'd80; 
32'd2672: dataIn2 = 32'd53; 
32'd2673: dataIn2 = 32'd38; 
32'd2674: dataIn2 = 32'd49; 
32'd2675: dataIn2 = 32'd55; 
32'd2676: dataIn2 = 32'd20; 
32'd2677: dataIn2 = 32'd13; 
32'd2678: dataIn2 = 32'd95; 
32'd2679: dataIn2 = 32'd64; 
32'd2680: dataIn2 = 32'd82; 
32'd2681: dataIn2 = 32'd39; 
32'd2682: dataIn2 = 32'd48; 
32'd2683: dataIn2 = 32'd66; 
32'd2684: dataIn2 = 32'd78; 
32'd2685: dataIn2 = 32'd92; 
32'd2686: dataIn2 = 32'd72; 
32'd2687: dataIn2 = 32'd49; 
32'd2688: dataIn2 = 32'd68; 
32'd2689: dataIn2 = 32'd73; 
32'd2690: dataIn2 = 32'd11; 
32'd2691: dataIn2 = 32'd47; 
32'd2692: dataIn2 = 32'd95; 
32'd2693: dataIn2 = 32'd83; 
32'd2694: dataIn2 = 32'd34; 
32'd2695: dataIn2 = 32'd85; 
32'd2696: dataIn2 = 32'd100; 
32'd2697: dataIn2 = 32'd45; 
32'd2698: dataIn2 = 32'd69; 
32'd2699: dataIn2 = 32'd12; 
32'd2700: dataIn2 = 32'd18; 
32'd2701: dataIn2 = 32'd94; 
32'd2702: dataIn2 = 32'd12; 
32'd2703: dataIn2 = 32'd33; 
32'd2704: dataIn2 = 32'd42; 
32'd2705: dataIn2 = 32'd3; 
32'd2706: dataIn2 = 32'd28; 
32'd2707: dataIn2 = 32'd21; 
32'd2708: dataIn2 = 32'd20; 
32'd2709: dataIn2 = 32'd93; 
32'd2710: dataIn2 = 32'd81; 
32'd2711: dataIn2 = 32'd5; 
32'd2712: dataIn2 = 32'd54; 
32'd2713: dataIn2 = 32'd32; 
32'd2714: dataIn2 = 32'd91; 
32'd2715: dataIn2 = 32'd69; 
32'd2716: dataIn2 = 32'd53; 
32'd2717: dataIn2 = 32'd68; 
32'd2718: dataIn2 = 32'd56; 
32'd2719: dataIn2 = 32'd81; 
32'd2720: dataIn2 = 32'd89; 
32'd2721: dataIn2 = 32'd88; 
32'd2722: dataIn2 = 32'd36; 
32'd2723: dataIn2 = 32'd87; 
32'd2724: dataIn2 = 32'd19; 
32'd2725: dataIn2 = 32'd38; 
32'd2726: dataIn2 = 32'd57; 
32'd2727: dataIn2 = 32'd68; 
32'd2728: dataIn2 = 32'd4; 
32'd2729: dataIn2 = 32'd73; 
32'd2730: dataIn2 = 32'd82; 
32'd2731: dataIn2 = 32'd84; 
32'd2732: dataIn2 = 32'd9; 
32'd2733: dataIn2 = 32'd11; 
32'd2734: dataIn2 = 32'd73; 
32'd2735: dataIn2 = 32'd38; 
32'd2736: dataIn2 = 32'd92; 
32'd2737: dataIn2 = 32'd80; 
32'd2738: dataIn2 = 32'd54; 
32'd2739: dataIn2 = 32'd32; 
32'd2740: dataIn2 = 32'd82; 
32'd2741: dataIn2 = 32'd39; 
32'd2742: dataIn2 = 32'd77; 
32'd2743: dataIn2 = 32'd2; 
32'd2744: dataIn2 = 32'd8; 
32'd2745: dataIn2 = 32'd37; 
32'd2746: dataIn2 = 32'd11; 
32'd2747: dataIn2 = 32'd83; 
32'd2748: dataIn2 = 32'd61; 
32'd2749: dataIn2 = 32'd49; 
32'd2750: dataIn2 = 32'd66; 
32'd2751: dataIn2 = 32'd30; 
32'd2752: dataIn2 = 32'd70; 
32'd2753: dataIn2 = 32'd50; 
32'd2754: dataIn2 = 32'd96; 
32'd2755: dataIn2 = 32'd37; 
32'd2756: dataIn2 = 32'd47; 
32'd2757: dataIn2 = 32'd11; 
32'd2758: dataIn2 = 32'd93; 
32'd2759: dataIn2 = 32'd58; 
32'd2760: dataIn2 = 32'd55; 
32'd2761: dataIn2 = 32'd1; 
32'd2762: dataIn2 = 32'd97; 
32'd2763: dataIn2 = 32'd73; 
32'd2764: dataIn2 = 32'd58; 
32'd2765: dataIn2 = 32'd97; 
32'd2766: dataIn2 = 32'd59; 
32'd2767: dataIn2 = 32'd2; 
32'd2768: dataIn2 = 32'd17; 
32'd2769: dataIn2 = 32'd21; 
32'd2770: dataIn2 = 32'd67; 
32'd2771: dataIn2 = 32'd81; 
32'd2772: dataIn2 = 32'd84; 
32'd2773: dataIn2 = 32'd78; 
32'd2774: dataIn2 = 32'd80; 
32'd2775: dataIn2 = 32'd27; 
32'd2776: dataIn2 = 32'd33; 
32'd2777: dataIn2 = 32'd68; 
32'd2778: dataIn2 = 32'd47; 
32'd2779: dataIn2 = 32'd37; 
32'd2780: dataIn2 = 32'd91; 
32'd2781: dataIn2 = 32'd18; 
32'd2782: dataIn2 = 32'd50; 
32'd2783: dataIn2 = 32'd36; 
32'd2784: dataIn2 = 32'd67; 
32'd2785: dataIn2 = 32'd55; 
32'd2786: dataIn2 = 32'd8; 
32'd2787: dataIn2 = 32'd0; 
32'd2788: dataIn2 = 32'd12; 
32'd2789: dataIn2 = 32'd30; 
32'd2790: dataIn2 = 32'd29; 
32'd2791: dataIn2 = 32'd37; 
32'd2792: dataIn2 = 32'd92; 
32'd2793: dataIn2 = 32'd74; 
32'd2794: dataIn2 = 32'd68; 
32'd2795: dataIn2 = 32'd95; 
32'd2796: dataIn2 = 32'd90; 
32'd2797: dataIn2 = 32'd6; 
32'd2798: dataIn2 = 32'd6; 
32'd2799: dataIn2 = 32'd54; 
32'd2800: dataIn2 = 32'd25; 
32'd2801: dataIn2 = 32'd1; 
32'd2802: dataIn2 = 32'd66; 
32'd2803: dataIn2 = 32'd76; 
32'd2804: dataIn2 = 32'd78; 
32'd2805: dataIn2 = 32'd53; 
32'd2806: dataIn2 = 32'd1; 
32'd2807: dataIn2 = 32'd93; 
32'd2808: dataIn2 = 32'd93; 
32'd2809: dataIn2 = 32'd2; 
32'd2810: dataIn2 = 32'd20; 
32'd2811: dataIn2 = 32'd10; 
32'd2812: dataIn2 = 32'd57; 
32'd2813: dataIn2 = 32'd88; 
32'd2814: dataIn2 = 32'd9; 
32'd2815: dataIn2 = 32'd53; 
32'd2816: dataIn2 = 32'd46; 
32'd2817: dataIn2 = 32'd8; 
32'd2818: dataIn2 = 32'd15; 
32'd2819: dataIn2 = 32'd99; 
32'd2820: dataIn2 = 32'd64; 
32'd2821: dataIn2 = 32'd28; 
32'd2822: dataIn2 = 32'd2; 
32'd2823: dataIn2 = 32'd65; 
32'd2824: dataIn2 = 32'd4; 
32'd2825: dataIn2 = 32'd61; 
32'd2826: dataIn2 = 32'd55; 
32'd2827: dataIn2 = 32'd26; 
32'd2828: dataIn2 = 32'd26; 
32'd2829: dataIn2 = 32'd65; 
32'd2830: dataIn2 = 32'd66; 
32'd2831: dataIn2 = 32'd66; 
32'd2832: dataIn2 = 32'd84; 
32'd2833: dataIn2 = 32'd100; 
32'd2834: dataIn2 = 32'd11; 
32'd2835: dataIn2 = 32'd15; 
32'd2836: dataIn2 = 32'd20; 
32'd2837: dataIn2 = 32'd80; 
32'd2838: dataIn2 = 32'd91; 
32'd2839: dataIn2 = 32'd31; 
32'd2840: dataIn2 = 32'd69; 
32'd2841: dataIn2 = 32'd56; 
32'd2842: dataIn2 = 32'd5; 
32'd2843: dataIn2 = 32'd73; 
32'd2844: dataIn2 = 32'd25; 
32'd2845: dataIn2 = 32'd7; 
32'd2846: dataIn2 = 32'd77; 
32'd2847: dataIn2 = 32'd78; 
32'd2848: dataIn2 = 32'd93; 
32'd2849: dataIn2 = 32'd68; 
32'd2850: dataIn2 = 32'd2; 
32'd2851: dataIn2 = 32'd45; 
32'd2852: dataIn2 = 32'd47; 
32'd2853: dataIn2 = 32'd83; 
32'd2854: dataIn2 = 32'd51; 
32'd2855: dataIn2 = 32'd62; 
32'd2856: dataIn2 = 32'd51; 
32'd2857: dataIn2 = 32'd84; 
32'd2858: dataIn2 = 32'd29; 
32'd2859: dataIn2 = 32'd66; 
32'd2860: dataIn2 = 32'd23; 
32'd2861: dataIn2 = 32'd63; 
32'd2862: dataIn2 = 32'd9; 
32'd2863: dataIn2 = 32'd97; 
32'd2864: dataIn2 = 32'd67; 
32'd2865: dataIn2 = 32'd21; 
32'd2866: dataIn2 = 32'd46; 
32'd2867: dataIn2 = 32'd21; 
32'd2868: dataIn2 = 32'd88; 
32'd2869: dataIn2 = 32'd84; 
32'd2870: dataIn2 = 32'd67; 
32'd2871: dataIn2 = 32'd6; 
32'd2872: dataIn2 = 32'd55; 
32'd2873: dataIn2 = 32'd37; 
32'd2874: dataIn2 = 32'd38; 
32'd2875: dataIn2 = 32'd84; 
32'd2876: dataIn2 = 32'd72; 
32'd2877: dataIn2 = 32'd88; 
32'd2878: dataIn2 = 32'd93; 
32'd2879: dataIn2 = 32'd3; 
32'd2880: dataIn2 = 32'd95; 
32'd2881: dataIn2 = 32'd1; 
32'd2882: dataIn2 = 32'd35; 
32'd2883: dataIn2 = 32'd3; 
32'd2884: dataIn2 = 32'd72; 
32'd2885: dataIn2 = 32'd54; 
32'd2886: dataIn2 = 32'd44; 
32'd2887: dataIn2 = 32'd36; 
32'd2888: dataIn2 = 32'd88; 
32'd2889: dataIn2 = 32'd86; 
32'd2890: dataIn2 = 32'd49; 
32'd2891: dataIn2 = 32'd77; 
32'd2892: dataIn2 = 32'd61; 
32'd2893: dataIn2 = 32'd76; 
32'd2894: dataIn2 = 32'd26; 
32'd2895: dataIn2 = 32'd0; 
32'd2896: dataIn2 = 32'd37; 
32'd2897: dataIn2 = 32'd75; 
32'd2898: dataIn2 = 32'd73; 
32'd2899: dataIn2 = 32'd4; 
32'd2900: dataIn2 = 32'd7; 
32'd2901: dataIn2 = 32'd10; 
32'd2902: dataIn2 = 32'd79; 
32'd2903: dataIn2 = 32'd36; 
32'd2904: dataIn2 = 32'd11; 
32'd2905: dataIn2 = 32'd35; 
32'd2906: dataIn2 = 32'd37; 
32'd2907: dataIn2 = 32'd65; 
32'd2908: dataIn2 = 32'd20; 
32'd2909: dataIn2 = 32'd22; 
32'd2910: dataIn2 = 32'd80; 
32'd2911: dataIn2 = 32'd75; 
32'd2912: dataIn2 = 32'd94; 
32'd2913: dataIn2 = 32'd57; 
32'd2914: dataIn2 = 32'd92; 
32'd2915: dataIn2 = 32'd28; 
32'd2916: dataIn2 = 32'd63; 
32'd2917: dataIn2 = 32'd66; 
32'd2918: dataIn2 = 32'd35; 
32'd2919: dataIn2 = 32'd12; 
32'd2920: dataIn2 = 32'd50; 
32'd2921: dataIn2 = 32'd80; 
32'd2922: dataIn2 = 32'd43; 
32'd2923: dataIn2 = 32'd45; 
32'd2924: dataIn2 = 32'd3; 
32'd2925: dataIn2 = 32'd13; 
32'd2926: dataIn2 = 32'd41; 
32'd2927: dataIn2 = 32'd35; 
32'd2928: dataIn2 = 32'd36; 
32'd2929: dataIn2 = 32'd83; 
32'd2930: dataIn2 = 32'd57; 
32'd2931: dataIn2 = 32'd55; 
32'd2932: dataIn2 = 32'd53; 
32'd2933: dataIn2 = 32'd59; 
32'd2934: dataIn2 = 32'd70; 
32'd2935: dataIn2 = 32'd100; 
32'd2936: dataIn2 = 32'd30; 
32'd2937: dataIn2 = 32'd97; 
32'd2938: dataIn2 = 32'd45; 
32'd2939: dataIn2 = 32'd88; 
32'd2940: dataIn2 = 32'd21; 
32'd2941: dataIn2 = 32'd78; 
32'd2942: dataIn2 = 32'd41; 
32'd2943: dataIn2 = 32'd68; 
32'd2944: dataIn2 = 32'd6; 
32'd2945: dataIn2 = 32'd13; 
32'd2946: dataIn2 = 32'd18; 
32'd2947: dataIn2 = 32'd23; 
32'd2948: dataIn2 = 32'd93; 
32'd2949: dataIn2 = 32'd9; 
32'd2950: dataIn2 = 32'd30; 
32'd2951: dataIn2 = 32'd64; 
32'd2952: dataIn2 = 32'd65; 
32'd2953: dataIn2 = 32'd25; 
32'd2954: dataIn2 = 32'd26; 
32'd2955: dataIn2 = 32'd94; 
32'd2956: dataIn2 = 32'd22; 
32'd2957: dataIn2 = 32'd88; 
32'd2958: dataIn2 = 32'd40; 
32'd2959: dataIn2 = 32'd7; 
32'd2960: dataIn2 = 32'd71; 
32'd2961: dataIn2 = 32'd54; 
32'd2962: dataIn2 = 32'd82; 
32'd2963: dataIn2 = 32'd75; 
32'd2964: dataIn2 = 32'd47; 
32'd2965: dataIn2 = 32'd67; 
32'd2966: dataIn2 = 32'd40; 
32'd2967: dataIn2 = 32'd99; 
32'd2968: dataIn2 = 32'd11; 
32'd2969: dataIn2 = 32'd85; 
32'd2970: dataIn2 = 32'd75; 
32'd2971: dataIn2 = 32'd28; 
32'd2972: dataIn2 = 32'd63; 
32'd2973: dataIn2 = 32'd72; 
32'd2974: dataIn2 = 32'd59; 
32'd2975: dataIn2 = 32'd97; 
32'd2976: dataIn2 = 32'd47; 
32'd2977: dataIn2 = 32'd81; 
32'd2978: dataIn2 = 32'd41; 
32'd2979: dataIn2 = 32'd7; 
32'd2980: dataIn2 = 32'd63; 
32'd2981: dataIn2 = 32'd79; 
32'd2982: dataIn2 = 32'd43; 
32'd2983: dataIn2 = 32'd54; 
32'd2984: dataIn2 = 32'd96; 
32'd2985: dataIn2 = 32'd71; 
32'd2986: dataIn2 = 32'd98; 
32'd2987: dataIn2 = 32'd59; 
32'd2988: dataIn2 = 32'd36; 
32'd2989: dataIn2 = 32'd20; 
32'd2990: dataIn2 = 32'd44; 
32'd2991: dataIn2 = 32'd59; 
32'd2992: dataIn2 = 32'd64; 
32'd2993: dataIn2 = 32'd55; 
32'd2994: dataIn2 = 32'd92; 
32'd2995: dataIn2 = 32'd28; 
32'd2996: dataIn2 = 32'd65; 
32'd2997: dataIn2 = 32'd46; 
32'd2998: dataIn2 = 32'd83; 
32'd2999: dataIn2 = 32'd45; 
32'd3000: dataIn2 = 32'd81; 
32'd3001: dataIn2 = 32'd69; 
32'd3002: dataIn2 = 32'd91; 
32'd3003: dataIn2 = 32'd70; 
32'd3004: dataIn2 = 32'd68; 
32'd3005: dataIn2 = 32'd81; 
32'd3006: dataIn2 = 32'd77; 
32'd3007: dataIn2 = 32'd96; 
32'd3008: dataIn2 = 32'd44; 
32'd3009: dataIn2 = 32'd85; 
32'd3010: dataIn2 = 32'd46; 
32'd3011: dataIn2 = 32'd43; 
32'd3012: dataIn2 = 32'd6; 
32'd3013: dataIn2 = 32'd58; 
32'd3014: dataIn2 = 32'd7; 
32'd3015: dataIn2 = 32'd93; 
32'd3016: dataIn2 = 32'd26; 
32'd3017: dataIn2 = 32'd43; 
32'd3018: dataIn2 = 32'd93; 
32'd3019: dataIn2 = 32'd14; 
32'd3020: dataIn2 = 32'd22; 
32'd3021: dataIn2 = 32'd5; 
32'd3022: dataIn2 = 32'd46; 
32'd3023: dataIn2 = 32'd87; 
32'd3024: dataIn2 = 32'd5; 
32'd3025: dataIn2 = 32'd53; 
32'd3026: dataIn2 = 32'd47; 
32'd3027: dataIn2 = 32'd15; 
32'd3028: dataIn2 = 32'd99; 
32'd3029: dataIn2 = 32'd65; 
32'd3030: dataIn2 = 32'd67; 
32'd3031: dataIn2 = 32'd0; 
32'd3032: dataIn2 = 32'd6; 
32'd3033: dataIn2 = 32'd2; 
32'd3034: dataIn2 = 32'd5; 
32'd3035: dataIn2 = 32'd6; 
32'd3036: dataIn2 = 32'd18; 
32'd3037: dataIn2 = 32'd63; 
32'd3038: dataIn2 = 32'd73; 
32'd3039: dataIn2 = 32'd6; 
32'd3040: dataIn2 = 32'd44; 
32'd3041: dataIn2 = 32'd34; 
32'd3042: dataIn2 = 32'd33; 
32'd3043: dataIn2 = 32'd68; 
32'd3044: dataIn2 = 32'd15; 
32'd3045: dataIn2 = 32'd23; 
32'd3046: dataIn2 = 32'd99; 
32'd3047: dataIn2 = 32'd34; 
32'd3048: dataIn2 = 32'd11; 
32'd3049: dataIn2 = 32'd25; 
32'd3050: dataIn2 = 32'd13; 
32'd3051: dataIn2 = 32'd30; 
32'd3052: dataIn2 = 32'd59; 
32'd3053: dataIn2 = 32'd63; 
32'd3054: dataIn2 = 32'd90; 
32'd3055: dataIn2 = 32'd85; 
32'd3056: dataIn2 = 32'd86; 
32'd3057: dataIn2 = 32'd57; 
32'd3058: dataIn2 = 32'd11; 
32'd3059: dataIn2 = 32'd84; 
32'd3060: dataIn2 = 32'd37; 
32'd3061: dataIn2 = 32'd60; 
32'd3062: dataIn2 = 32'd17; 
32'd3063: dataIn2 = 32'd72; 
32'd3064: dataIn2 = 32'd2; 
32'd3065: dataIn2 = 32'd34; 
32'd3066: dataIn2 = 32'd31; 
32'd3067: dataIn2 = 32'd31; 
32'd3068: dataIn2 = 32'd8; 
32'd3069: dataIn2 = 32'd11; 
32'd3070: dataIn2 = 32'd97; 
32'd3071: dataIn2 = 32'd0; 
32'd3072: dataIn2 = 32'd86; 
32'd3073: dataIn2 = 32'd83; 
32'd3074: dataIn2 = 32'd17; 
32'd3075: dataIn2 = 32'd55; 
32'd3076: dataIn2 = 32'd19; 
32'd3077: dataIn2 = 32'd77; 
32'd3078: dataIn2 = 32'd43; 
32'd3079: dataIn2 = 32'd5; 
32'd3080: dataIn2 = 32'd98; 
32'd3081: dataIn2 = 32'd14; 
32'd3082: dataIn2 = 32'd11; 
32'd3083: dataIn2 = 32'd18; 
32'd3084: dataIn2 = 32'd80; 
32'd3085: dataIn2 = 32'd65; 
32'd3086: dataIn2 = 32'd48; 
32'd3087: dataIn2 = 32'd96; 
32'd3088: dataIn2 = 32'd50; 
32'd3089: dataIn2 = 32'd4; 
32'd3090: dataIn2 = 32'd9; 
32'd3091: dataIn2 = 32'd7; 
32'd3092: dataIn2 = 32'd28; 
32'd3093: dataIn2 = 32'd9; 
32'd3094: dataIn2 = 32'd100; 
32'd3095: dataIn2 = 32'd96; 
32'd3096: dataIn2 = 32'd73; 
32'd3097: dataIn2 = 32'd72; 
32'd3098: dataIn2 = 32'd40; 
32'd3099: dataIn2 = 32'd23; 
32'd3100: dataIn2 = 32'd68; 
32'd3101: dataIn2 = 32'd49; 
32'd3102: dataIn2 = 32'd89; 
32'd3103: dataIn2 = 32'd11; 
32'd3104: dataIn2 = 32'd7; 
32'd3105: dataIn2 = 32'd49; 
32'd3106: dataIn2 = 32'd92; 
32'd3107: dataIn2 = 32'd13; 
32'd3108: dataIn2 = 32'd70; 
32'd3109: dataIn2 = 32'd71; 
32'd3110: dataIn2 = 32'd11; 
32'd3111: dataIn2 = 32'd11; 
32'd3112: dataIn2 = 32'd6; 
32'd3113: dataIn2 = 32'd12; 
32'd3114: dataIn2 = 32'd80; 
32'd3115: dataIn2 = 32'd19; 
32'd3116: dataIn2 = 32'd98; 
32'd3117: dataIn2 = 32'd52; 
32'd3118: dataIn2 = 32'd18; 
32'd3119: dataIn2 = 32'd84; 
32'd3120: dataIn2 = 32'd27; 
32'd3121: dataIn2 = 32'd42; 
32'd3122: dataIn2 = 32'd15; 
32'd3123: dataIn2 = 32'd2; 
32'd3124: dataIn2 = 32'd80; 
32'd3125: dataIn2 = 32'd10; 
32'd3126: dataIn2 = 32'd6; 
32'd3127: dataIn2 = 32'd66; 
32'd3128: dataIn2 = 32'd69; 
32'd3129: dataIn2 = 32'd18; 
32'd3130: dataIn2 = 32'd25; 
32'd3131: dataIn2 = 32'd34; 
32'd3132: dataIn2 = 32'd55; 
32'd3133: dataIn2 = 32'd50; 
32'd3134: dataIn2 = 32'd13; 
32'd3135: dataIn2 = 32'd77; 
32'd3136: dataIn2 = 32'd58; 
32'd3137: dataIn2 = 32'd79; 
32'd3138: dataIn2 = 32'd91; 
32'd3139: dataIn2 = 32'd29; 
32'd3140: dataIn2 = 32'd73; 
32'd3141: dataIn2 = 32'd78; 
32'd3142: dataIn2 = 32'd98; 
32'd3143: dataIn2 = 32'd73; 
32'd3144: dataIn2 = 32'd8; 
32'd3145: dataIn2 = 32'd79; 
32'd3146: dataIn2 = 32'd89; 
32'd3147: dataIn2 = 32'd53; 
32'd3148: dataIn2 = 32'd94; 
32'd3149: dataIn2 = 32'd99; 
32'd3150: dataIn2 = 32'd31; 
32'd3151: dataIn2 = 32'd4; 
32'd3152: dataIn2 = 32'd45; 
32'd3153: dataIn2 = 32'd84; 
32'd3154: dataIn2 = 32'd37; 
32'd3155: dataIn2 = 32'd91; 
32'd3156: dataIn2 = 32'd42; 
32'd3157: dataIn2 = 32'd10; 
32'd3158: dataIn2 = 32'd68; 
32'd3159: dataIn2 = 32'd50; 
32'd3160: dataIn2 = 32'd87; 
32'd3161: dataIn2 = 32'd87; 
32'd3162: dataIn2 = 32'd6; 
32'd3163: dataIn2 = 32'd11; 
32'd3164: dataIn2 = 32'd89; 
32'd3165: dataIn2 = 32'd64; 
32'd3166: dataIn2 = 32'd88; 
32'd3167: dataIn2 = 32'd69; 
32'd3168: dataIn2 = 32'd93; 
32'd3169: dataIn2 = 32'd41; 
32'd3170: dataIn2 = 32'd0; 
32'd3171: dataIn2 = 32'd2; 
32'd3172: dataIn2 = 32'd22; 
32'd3173: dataIn2 = 32'd71; 
32'd3174: dataIn2 = 32'd37; 
32'd3175: dataIn2 = 32'd79; 
32'd3176: dataIn2 = 32'd9; 
32'd3177: dataIn2 = 32'd39; 
32'd3178: dataIn2 = 32'd100; 
32'd3179: dataIn2 = 32'd2; 
32'd3180: dataIn2 = 32'd25; 
32'd3181: dataIn2 = 32'd81; 
32'd3182: dataIn2 = 32'd17; 
32'd3183: dataIn2 = 32'd79; 
32'd3184: dataIn2 = 32'd89; 
32'd3185: dataIn2 = 32'd94; 
32'd3186: dataIn2 = 32'd2; 
32'd3187: dataIn2 = 32'd78; 
32'd3188: dataIn2 = 32'd2; 
32'd3189: dataIn2 = 32'd5; 
32'd3190: dataIn2 = 32'd83; 
32'd3191: dataIn2 = 32'd72; 
32'd3192: dataIn2 = 32'd31; 
32'd3193: dataIn2 = 32'd13; 
32'd3194: dataIn2 = 32'd100; 
32'd3195: dataIn2 = 32'd6; 
32'd3196: dataIn2 = 32'd100; 
32'd3197: dataIn2 = 32'd52; 
32'd3198: dataIn2 = 32'd30; 
32'd3199: dataIn2 = 32'd9; 
32'd3200: dataIn2 = 32'd99; 
32'd3201: dataIn2 = 32'd59; 
32'd3202: dataIn2 = 32'd77; 
32'd3203: dataIn2 = 32'd72; 
32'd3204: dataIn2 = 32'd25; 
32'd3205: dataIn2 = 32'd38; 
32'd3206: dataIn2 = 32'd55; 
32'd3207: dataIn2 = 32'd72; 
32'd3208: dataIn2 = 32'd89; 
32'd3209: dataIn2 = 32'd78; 
32'd3210: dataIn2 = 32'd13; 
32'd3211: dataIn2 = 32'd72; 
32'd3212: dataIn2 = 32'd42; 
32'd3213: dataIn2 = 32'd88; 
32'd3214: dataIn2 = 32'd63; 
32'd3215: dataIn2 = 32'd80; 
32'd3216: dataIn2 = 32'd64; 
32'd3217: dataIn2 = 32'd97; 
32'd3218: dataIn2 = 32'd60; 
32'd3219: dataIn2 = 32'd0; 
32'd3220: dataIn2 = 32'd38; 
32'd3221: dataIn2 = 32'd51; 
32'd3222: dataIn2 = 32'd94; 
32'd3223: dataIn2 = 32'd66; 
32'd3224: dataIn2 = 32'd98; 
32'd3225: dataIn2 = 32'd34; 
32'd3226: dataIn2 = 32'd90; 
32'd3227: dataIn2 = 32'd67; 
32'd3228: dataIn2 = 32'd13; 
32'd3229: dataIn2 = 32'd16; 
32'd3230: dataIn2 = 32'd70; 
32'd3231: dataIn2 = 32'd64; 
32'd3232: dataIn2 = 32'd55; 
32'd3233: dataIn2 = 32'd45; 
32'd3234: dataIn2 = 32'd2; 
32'd3235: dataIn2 = 32'd6; 
32'd3236: dataIn2 = 32'd89; 
32'd3237: dataIn2 = 32'd11; 
32'd3238: dataIn2 = 32'd94; 
32'd3239: dataIn2 = 32'd9; 
32'd3240: dataIn2 = 32'd60; 
32'd3241: dataIn2 = 32'd97; 
32'd3242: dataIn2 = 32'd47; 
32'd3243: dataIn2 = 32'd3; 
32'd3244: dataIn2 = 32'd8; 
32'd3245: dataIn2 = 32'd27; 
32'd3246: dataIn2 = 32'd79; 
32'd3247: dataIn2 = 32'd51; 
32'd3248: dataIn2 = 32'd29; 
32'd3249: dataIn2 = 32'd14; 
32'd3250: dataIn2 = 32'd15; 
32'd3251: dataIn2 = 32'd81; 
32'd3252: dataIn2 = 32'd54; 
32'd3253: dataIn2 = 32'd5; 
32'd3254: dataIn2 = 32'd79; 
32'd3255: dataIn2 = 32'd51; 
32'd3256: dataIn2 = 32'd81; 
32'd3257: dataIn2 = 32'd57; 
32'd3258: dataIn2 = 32'd100; 
32'd3259: dataIn2 = 32'd93; 
32'd3260: dataIn2 = 32'd9; 
32'd3261: dataIn2 = 32'd56; 
32'd3262: dataIn2 = 32'd64; 
32'd3263: dataIn2 = 32'd33; 
32'd3264: dataIn2 = 32'd90; 
32'd3265: dataIn2 = 32'd61; 
32'd3266: dataIn2 = 32'd63; 
32'd3267: dataIn2 = 32'd100; 
32'd3268: dataIn2 = 32'd17; 
32'd3269: dataIn2 = 32'd71; 
32'd3270: dataIn2 = 32'd84; 
32'd3271: dataIn2 = 32'd86; 
32'd3272: dataIn2 = 32'd10; 
32'd3273: dataIn2 = 32'd7; 
32'd3274: dataIn2 = 32'd10; 
32'd3275: dataIn2 = 32'd34; 
32'd3276: dataIn2 = 32'd45; 
32'd3277: dataIn2 = 32'd4; 
32'd3278: dataIn2 = 32'd97; 
32'd3279: dataIn2 = 32'd91; 
32'd3280: dataIn2 = 32'd23; 
32'd3281: dataIn2 = 32'd48; 
32'd3282: dataIn2 = 32'd5; 
32'd3283: dataIn2 = 32'd40; 
32'd3284: dataIn2 = 32'd9; 
32'd3285: dataIn2 = 32'd100; 
32'd3286: dataIn2 = 32'd1; 
32'd3287: dataIn2 = 32'd26; 
32'd3288: dataIn2 = 32'd39; 
32'd3289: dataIn2 = 32'd61; 
32'd3290: dataIn2 = 32'd85; 
32'd3291: dataIn2 = 32'd60; 
32'd3292: dataIn2 = 32'd75; 
32'd3293: dataIn2 = 32'd25; 
32'd3294: dataIn2 = 32'd42; 
32'd3295: dataIn2 = 32'd80; 
32'd3296: dataIn2 = 32'd54; 
32'd3297: dataIn2 = 32'd17; 
32'd3298: dataIn2 = 32'd23; 
32'd3299: dataIn2 = 32'd62; 
32'd3300: dataIn2 = 32'd8; 
32'd3301: dataIn2 = 32'd60; 
32'd3302: dataIn2 = 32'd56; 
32'd3303: dataIn2 = 32'd64; 
32'd3304: dataIn2 = 32'd12; 
32'd3305: dataIn2 = 32'd79; 
32'd3306: dataIn2 = 32'd40; 
32'd3307: dataIn2 = 32'd23; 
32'd3308: dataIn2 = 32'd64; 
32'd3309: dataIn2 = 32'd58; 
32'd3310: dataIn2 = 32'd90; 
32'd3311: dataIn2 = 32'd73; 
32'd3312: dataIn2 = 32'd7; 
32'd3313: dataIn2 = 32'd93; 
32'd3314: dataIn2 = 32'd32; 
32'd3315: dataIn2 = 32'd81; 
32'd3316: dataIn2 = 32'd4; 
32'd3317: dataIn2 = 32'd85; 
32'd3318: dataIn2 = 32'd93; 
32'd3319: dataIn2 = 32'd15; 
32'd3320: dataIn2 = 32'd91; 
32'd3321: dataIn2 = 32'd90; 
32'd3322: dataIn2 = 32'd96; 
32'd3323: dataIn2 = 32'd71; 
32'd3324: dataIn2 = 32'd7; 
32'd3325: dataIn2 = 32'd23; 
32'd3326: dataIn2 = 32'd29; 
32'd3327: dataIn2 = 32'd36; 
32'd3328: dataIn2 = 32'd62; 
32'd3329: dataIn2 = 32'd80; 
32'd3330: dataIn2 = 32'd57; 
32'd3331: dataIn2 = 32'd9; 
32'd3332: dataIn2 = 32'd92; 
32'd3333: dataIn2 = 32'd26; 
32'd3334: dataIn2 = 32'd46; 
32'd3335: dataIn2 = 32'd28; 
32'd3336: dataIn2 = 32'd32; 
32'd3337: dataIn2 = 32'd23; 
32'd3338: dataIn2 = 32'd44; 
32'd3339: dataIn2 = 32'd3; 
32'd3340: dataIn2 = 32'd86; 
32'd3341: dataIn2 = 32'd48; 
32'd3342: dataIn2 = 32'd43; 
32'd3343: dataIn2 = 32'd59; 
32'd3344: dataIn2 = 32'd47; 
32'd3345: dataIn2 = 32'd52; 
32'd3346: dataIn2 = 32'd23; 
32'd3347: dataIn2 = 32'd82; 
32'd3348: dataIn2 = 32'd98; 
32'd3349: dataIn2 = 32'd22; 
32'd3350: dataIn2 = 32'd67; 
32'd3351: dataIn2 = 32'd55; 
32'd3352: dataIn2 = 32'd51; 
32'd3353: dataIn2 = 32'd19; 
32'd3354: dataIn2 = 32'd47; 
32'd3355: dataIn2 = 32'd21; 
32'd3356: dataIn2 = 32'd3; 
32'd3357: dataIn2 = 32'd84; 
32'd3358: dataIn2 = 32'd58; 
32'd3359: dataIn2 = 32'd59; 
32'd3360: dataIn2 = 32'd25; 
32'd3361: dataIn2 = 32'd82; 
32'd3362: dataIn2 = 32'd94; 
32'd3363: dataIn2 = 32'd4; 
32'd3364: dataIn2 = 32'd95; 
32'd3365: dataIn2 = 32'd48; 
32'd3366: dataIn2 = 32'd61; 
32'd3367: dataIn2 = 32'd15; 
32'd3368: dataIn2 = 32'd74; 
32'd3369: dataIn2 = 32'd87; 
32'd3370: dataIn2 = 32'd99; 
32'd3371: dataIn2 = 32'd12; 
32'd3372: dataIn2 = 32'd100; 
32'd3373: dataIn2 = 32'd25; 
32'd3374: dataIn2 = 32'd3; 
32'd3375: dataIn2 = 32'd65; 
32'd3376: dataIn2 = 32'd21; 
32'd3377: dataIn2 = 32'd12; 
32'd3378: dataIn2 = 32'd39; 
32'd3379: dataIn2 = 32'd70; 
32'd3380: dataIn2 = 32'd37; 
32'd3381: dataIn2 = 32'd32; 
32'd3382: dataIn2 = 32'd5; 
32'd3383: dataIn2 = 32'd21; 
32'd3384: dataIn2 = 32'd68; 
32'd3385: dataIn2 = 32'd81; 
32'd3386: dataIn2 = 32'd61; 
32'd3387: dataIn2 = 32'd28; 
32'd3388: dataIn2 = 32'd83; 
32'd3389: dataIn2 = 32'd84; 
32'd3390: dataIn2 = 32'd16; 
32'd3391: dataIn2 = 32'd60; 
32'd3392: dataIn2 = 32'd69; 
32'd3393: dataIn2 = 32'd29; 
32'd3394: dataIn2 = 32'd8; 
32'd3395: dataIn2 = 32'd53; 
32'd3396: dataIn2 = 32'd25; 
32'd3397: dataIn2 = 32'd45; 
32'd3398: dataIn2 = 32'd23; 
32'd3399: dataIn2 = 32'd68; 
32'd3400: dataIn2 = 32'd97; 
32'd3401: dataIn2 = 32'd1; 
32'd3402: dataIn2 = 32'd24; 
32'd3403: dataIn2 = 32'd32; 
32'd3404: dataIn2 = 32'd0; 
32'd3405: dataIn2 = 32'd69; 
32'd3406: dataIn2 = 32'd63; 
32'd3407: dataIn2 = 32'd90; 
32'd3408: dataIn2 = 32'd83; 
32'd3409: dataIn2 = 32'd76; 
32'd3410: dataIn2 = 32'd55; 
32'd3411: dataIn2 = 32'd57; 
32'd3412: dataIn2 = 32'd75; 
32'd3413: dataIn2 = 32'd69; 
32'd3414: dataIn2 = 32'd28; 
32'd3415: dataIn2 = 32'd34; 
32'd3416: dataIn2 = 32'd52; 
32'd3417: dataIn2 = 32'd58; 
32'd3418: dataIn2 = 32'd35; 
32'd3419: dataIn2 = 32'd92; 
32'd3420: dataIn2 = 32'd38; 
32'd3421: dataIn2 = 32'd11; 
32'd3422: dataIn2 = 32'd93; 
32'd3423: dataIn2 = 32'd9; 
32'd3424: dataIn2 = 32'd9; 
32'd3425: dataIn2 = 32'd9; 
32'd3426: dataIn2 = 32'd59; 
32'd3427: dataIn2 = 32'd62; 
32'd3428: dataIn2 = 32'd91; 
32'd3429: dataIn2 = 32'd82; 
32'd3430: dataIn2 = 32'd48; 
32'd3431: dataIn2 = 32'd51; 
32'd3432: dataIn2 = 32'd91; 
32'd3433: dataIn2 = 32'd100; 
32'd3434: dataIn2 = 32'd95; 
32'd3435: dataIn2 = 32'd1; 
32'd3436: dataIn2 = 32'd3; 
32'd3437: dataIn2 = 32'd86; 
32'd3438: dataIn2 = 32'd42; 
32'd3439: dataIn2 = 32'd7; 
32'd3440: dataIn2 = 32'd45; 
32'd3441: dataIn2 = 32'd89; 
32'd3442: dataIn2 = 32'd96; 
32'd3443: dataIn2 = 32'd30; 
32'd3444: dataIn2 = 32'd99; 
32'd3445: dataIn2 = 32'd17; 
32'd3446: dataIn2 = 32'd91; 
32'd3447: dataIn2 = 32'd11; 
32'd3448: dataIn2 = 32'd14; 
32'd3449: dataIn2 = 32'd15; 
32'd3450: dataIn2 = 32'd50; 
32'd3451: dataIn2 = 32'd3; 
32'd3452: dataIn2 = 32'd59; 
32'd3453: dataIn2 = 32'd79; 
32'd3454: dataIn2 = 32'd70; 
32'd3455: dataIn2 = 32'd45; 
32'd3456: dataIn2 = 32'd14; 
32'd3457: dataIn2 = 32'd21; 
32'd3458: dataIn2 = 32'd1; 
32'd3459: dataIn2 = 32'd10; 
32'd3460: dataIn2 = 32'd3; 
32'd3461: dataIn2 = 32'd65; 
32'd3462: dataIn2 = 32'd6; 
32'd3463: dataIn2 = 32'd12; 
32'd3464: dataIn2 = 32'd10; 
32'd3465: dataIn2 = 32'd57; 
32'd3466: dataIn2 = 32'd66; 
32'd3467: dataIn2 = 32'd29; 
32'd3468: dataIn2 = 32'd30; 
32'd3469: dataIn2 = 32'd91; 
32'd3470: dataIn2 = 32'd19; 
32'd3471: dataIn2 = 32'd62; 
32'd3472: dataIn2 = 32'd66; 
32'd3473: dataIn2 = 32'd57; 
32'd3474: dataIn2 = 32'd74; 
32'd3475: dataIn2 = 32'd75; 
32'd3476: dataIn2 = 32'd69; 
32'd3477: dataIn2 = 32'd60; 
32'd3478: dataIn2 = 32'd93; 
32'd3479: dataIn2 = 32'd64; 
32'd3480: dataIn2 = 32'd46; 
32'd3481: dataIn2 = 32'd35; 
32'd3482: dataIn2 = 32'd42; 
32'd3483: dataIn2 = 32'd94; 
32'd3484: dataIn2 = 32'd79; 
32'd3485: dataIn2 = 32'd40; 
32'd3486: dataIn2 = 32'd53; 
32'd3487: dataIn2 = 32'd98; 
32'd3488: dataIn2 = 32'd0; 
32'd3489: dataIn2 = 32'd75; 
32'd3490: dataIn2 = 32'd5; 
32'd3491: dataIn2 = 32'd87; 
32'd3492: dataIn2 = 32'd20; 
32'd3493: dataIn2 = 32'd43; 
32'd3494: dataIn2 = 32'd94; 
32'd3495: dataIn2 = 32'd44; 
32'd3496: dataIn2 = 32'd69; 
32'd3497: dataIn2 = 32'd45; 
32'd3498: dataIn2 = 32'd95; 
32'd3499: dataIn2 = 32'd73; 
32'd3500: dataIn2 = 32'd60; 
32'd3501: dataIn2 = 32'd37; 
32'd3502: dataIn2 = 32'd84; 
32'd3503: dataIn2 = 32'd57; 
32'd3504: dataIn2 = 32'd93; 
32'd3505: dataIn2 = 32'd92; 
32'd3506: dataIn2 = 32'd46; 
32'd3507: dataIn2 = 32'd15; 
32'd3508: dataIn2 = 32'd67; 
32'd3509: dataIn2 = 32'd85; 
32'd3510: dataIn2 = 32'd56; 
32'd3511: dataIn2 = 32'd59; 
32'd3512: dataIn2 = 32'd9; 
32'd3513: dataIn2 = 32'd39; 
32'd3514: dataIn2 = 32'd21; 
32'd3515: dataIn2 = 32'd85; 
32'd3516: dataIn2 = 32'd16; 
32'd3517: dataIn2 = 32'd47; 
32'd3518: dataIn2 = 32'd99; 
32'd3519: dataIn2 = 32'd76; 
32'd3520: dataIn2 = 32'd81; 
32'd3521: dataIn2 = 32'd65; 
32'd3522: dataIn2 = 32'd59; 
32'd3523: dataIn2 = 32'd50; 
32'd3524: dataIn2 = 32'd48; 
32'd3525: dataIn2 = 32'd29; 
32'd3526: dataIn2 = 32'd61; 
32'd3527: dataIn2 = 32'd71; 
32'd3528: dataIn2 = 32'd85; 
32'd3529: dataIn2 = 32'd60; 
32'd3530: dataIn2 = 32'd98; 
32'd3531: dataIn2 = 32'd53; 
32'd3532: dataIn2 = 32'd79; 
32'd3533: dataIn2 = 32'd6; 
32'd3534: dataIn2 = 32'd85; 
32'd3535: dataIn2 = 32'd76; 
32'd3536: dataIn2 = 32'd53; 
32'd3537: dataIn2 = 32'd74; 
32'd3538: dataIn2 = 32'd71; 
32'd3539: dataIn2 = 32'd28; 
32'd3540: dataIn2 = 32'd27; 
32'd3541: dataIn2 = 32'd90; 
32'd3542: dataIn2 = 32'd16; 
32'd3543: dataIn2 = 32'd95; 
32'd3544: dataIn2 = 32'd18; 
32'd3545: dataIn2 = 32'd25; 
32'd3546: dataIn2 = 32'd85; 
32'd3547: dataIn2 = 32'd99; 
32'd3548: dataIn2 = 32'd37; 
32'd3549: dataIn2 = 32'd93; 
32'd3550: dataIn2 = 32'd58; 
32'd3551: dataIn2 = 32'd9; 
32'd3552: dataIn2 = 32'd50; 
32'd3553: dataIn2 = 32'd66; 
32'd3554: dataIn2 = 32'd53; 
32'd3555: dataIn2 = 32'd56; 
32'd3556: dataIn2 = 32'd51; 
32'd3557: dataIn2 = 32'd91; 
32'd3558: dataIn2 = 32'd44; 
32'd3559: dataIn2 = 32'd0; 
32'd3560: dataIn2 = 32'd46; 
32'd3561: dataIn2 = 32'd76; 
32'd3562: dataIn2 = 32'd73; 
32'd3563: dataIn2 = 32'd76; 
32'd3564: dataIn2 = 32'd12; 
32'd3565: dataIn2 = 32'd3; 
32'd3566: dataIn2 = 32'd95; 
32'd3567: dataIn2 = 32'd59; 
32'd3568: dataIn2 = 32'd36; 
32'd3569: dataIn2 = 32'd66; 
32'd3570: dataIn2 = 32'd32; 
32'd3571: dataIn2 = 32'd21; 
32'd3572: dataIn2 = 32'd37; 
32'd3573: dataIn2 = 32'd11; 
32'd3574: dataIn2 = 32'd23; 
32'd3575: dataIn2 = 32'd86; 
32'd3576: dataIn2 = 32'd39; 
32'd3577: dataIn2 = 32'd64; 
32'd3578: dataIn2 = 32'd44; 
32'd3579: dataIn2 = 32'd41; 
32'd3580: dataIn2 = 32'd73; 
32'd3581: dataIn2 = 32'd71; 
32'd3582: dataIn2 = 32'd0; 
32'd3583: dataIn2 = 32'd19; 
32'd3584: dataIn2 = 32'd55; 
32'd3585: dataIn2 = 32'd76; 
32'd3586: dataIn2 = 32'd87; 
32'd3587: dataIn2 = 32'd51; 
32'd3588: dataIn2 = 32'd51; 
32'd3589: dataIn2 = 32'd40; 
32'd3590: dataIn2 = 32'd12; 
32'd3591: dataIn2 = 32'd19; 
32'd3592: dataIn2 = 32'd31; 
32'd3593: dataIn2 = 32'd83; 
32'd3594: dataIn2 = 32'd85; 
32'd3595: dataIn2 = 32'd57; 
32'd3596: dataIn2 = 32'd82; 
32'd3597: dataIn2 = 32'd28; 
32'd3598: dataIn2 = 32'd78; 
32'd3599: dataIn2 = 32'd100; 
32'd3600: dataIn2 = 32'd100; 
32'd3601: dataIn2 = 32'd97; 
32'd3602: dataIn2 = 32'd51; 
32'd3603: dataIn2 = 32'd21; 
32'd3604: dataIn2 = 32'd9; 
32'd3605: dataIn2 = 32'd76; 
32'd3606: dataIn2 = 32'd93; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_64_20.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
