//32x32 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 410 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd170 ; 
  wdata_col_base = 32'd5800 ; 
  row_base = 32'd62100 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #8380; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd62100: dataIn1 = 32'd0
; 
32'd62101: dataIn1 = 32'd17
; 
32'd62102: dataIn1 = 32'd27
; 
32'd62103: dataIn1 = 32'd36
; 
32'd62104: dataIn1 = 32'd47
; 
32'd62105: dataIn1 = 32'd58
; 
32'd62106: dataIn1 = 32'd70
; 
32'd62107: dataIn1 = 32'd83
; 
32'd62108: dataIn1 = 32'd100
; 
32'd62109: dataIn1 = 32'd111
; 
32'd62110: dataIn1 = 32'd122
; 
32'd62111: dataIn1 = 32'd133
; 
32'd62112: dataIn1 = 32'd149
; 
32'd62113: dataIn1 = 32'd159
; 
32'd62114: dataIn1 = 32'd177
; 
32'd62115: dataIn1 = 32'd189
; 
32'd62116: dataIn1 = 32'd200
; 
32'd62117: dataIn1 = 32'd207
; 
32'd62118: dataIn1 = 32'd220
; 
32'd62119: dataIn1 = 32'd233
; 
32'd62120: dataIn1 = 32'd244
; 
32'd62121: dataIn1 = 32'd257
; 
32'd62122: dataIn1 = 32'd265
; 
32'd62123: dataIn1 = 32'd278
; 
32'd62124: dataIn1 = 32'd292
; 
32'd62125: dataIn1 = 32'd302
; 
32'd62126: dataIn1 = 32'd311
; 
32'd62127: dataIn1 = 32'd317
; 
32'd62128: dataIn1 = 32'd332
; 
32'd62129: dataIn1 = 32'd346
; 
32'd62130: dataIn1 = 32'd360
; 
32'd62131: dataIn1 = 32'd375
; 
32'd62132: dataIn1 = 32'd385
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd5800: dataIn1 = 32'd0
; 
32'd5801: dataIn1 = 32'd17
; 
32'd5802: dataIn1 = 32'd27
; 
32'd5803: dataIn1 = 32'd36
; 
32'd5804: dataIn1 = 32'd47
; 
32'd5805: dataIn1 = 32'd58
; 
32'd5806: dataIn1 = 32'd70
; 
32'd5807: dataIn1 = 32'd83
; 
32'd5808: dataIn1 = 32'd100
; 
32'd5809: dataIn1 = 32'd111
; 
32'd5810: dataIn1 = 32'd122
; 
32'd5811: dataIn1 = 32'd133
; 
32'd5812: dataIn1 = 32'd149
; 
32'd5813: dataIn1 = 32'd159
; 
32'd5814: dataIn1 = 32'd177
; 
32'd5815: dataIn1 = 32'd189
; 
32'd5816: dataIn1 = 32'd200
; 
32'd5817: dataIn1 = 32'd207
; 
32'd5818: dataIn1 = 32'd220
; 
32'd5819: dataIn1 = 32'd233
; 
32'd5820: dataIn1 = 32'd244
; 
32'd5821: dataIn1 = 32'd257
; 
32'd5822: dataIn1 = 32'd265
; 
32'd5823: dataIn1 = 32'd278
; 
32'd5824: dataIn1 = 32'd292
; 
32'd5825: dataIn1 = 32'd302
; 
32'd5826: dataIn1 = 32'd311
; 
32'd5827: dataIn1 = 32'd317
; 
32'd5828: dataIn1 = 32'd332
; 
32'd5829: dataIn1 = 32'd346
; 
32'd5830: dataIn1 = 32'd360
; 
32'd5831: dataIn1 = 32'd375
; 
32'd5832: dataIn1 = 32'd385
; 
32'd5833: dataIn1 = 32'd3
; 
32'd5834: dataIn1 = 32'd4
; 
32'd5835: dataIn1 = 32'd5
; 
32'd5836: dataIn1 = 32'd6
; 
32'd5837: dataIn1 = 32'd8
; 
32'd5838: dataIn1 = 32'd10
; 
32'd5839: dataIn1 = 32'd12
; 
32'd5840: dataIn1 = 32'd13
; 
32'd5841: dataIn1 = 32'd15
; 
32'd5842: dataIn1 = 32'd17
; 
32'd5843: dataIn1 = 32'd19
; 
32'd5844: dataIn1 = 32'd20
; 
32'd5845: dataIn1 = 32'd21
; 
32'd5846: dataIn1 = 32'd23
; 
32'd5847: dataIn1 = 32'd26
; 
32'd5848: dataIn1 = 32'd27
; 
32'd5849: dataIn1 = 32'd30
; 
32'd5850: dataIn1 = 32'd0
; 
32'd5851: dataIn1 = 32'd4
; 
32'd5852: dataIn1 = 32'd5
; 
32'd5853: dataIn1 = 32'd6
; 
32'd5854: dataIn1 = 32'd11
; 
32'd5855: dataIn1 = 32'd12
; 
32'd5856: dataIn1 = 32'd19
; 
32'd5857: dataIn1 = 32'd24
; 
32'd5858: dataIn1 = 32'd28
; 
32'd5859: dataIn1 = 32'd29
; 
32'd5860: dataIn1 = 32'd1
; 
32'd5861: dataIn1 = 32'd6
; 
32'd5862: dataIn1 = 32'd9
; 
32'd5863: dataIn1 = 32'd18
; 
32'd5864: dataIn1 = 32'd19
; 
32'd5865: dataIn1 = 32'd20
; 
32'd5866: dataIn1 = 32'd21
; 
32'd5867: dataIn1 = 32'd29
; 
32'd5868: dataIn1 = 32'd31
; 
32'd5869: dataIn1 = 32'd5
; 
32'd5870: dataIn1 = 32'd6
; 
32'd5871: dataIn1 = 32'd8
; 
32'd5872: dataIn1 = 32'd9
; 
32'd5873: dataIn1 = 32'd11
; 
32'd5874: dataIn1 = 32'd12
; 
32'd5875: dataIn1 = 32'd14
; 
32'd5876: dataIn1 = 32'd19
; 
32'd5877: dataIn1 = 32'd22
; 
32'd5878: dataIn1 = 32'd26
; 
32'd5879: dataIn1 = 32'd27
; 
32'd5880: dataIn1 = 32'd4
; 
32'd5881: dataIn1 = 32'd5
; 
32'd5882: dataIn1 = 32'd6
; 
32'd5883: dataIn1 = 32'd10
; 
32'd5884: dataIn1 = 32'd14
; 
32'd5885: dataIn1 = 32'd17
; 
32'd5886: dataIn1 = 32'd18
; 
32'd5887: dataIn1 = 32'd20
; 
32'd5888: dataIn1 = 32'd24
; 
32'd5889: dataIn1 = 32'd27
; 
32'd5890: dataIn1 = 32'd30
; 
32'd5891: dataIn1 = 32'd4
; 
32'd5892: dataIn1 = 32'd5
; 
32'd5893: dataIn1 = 32'd8
; 
32'd5894: dataIn1 = 32'd13
; 
32'd5895: dataIn1 = 32'd15
; 
32'd5896: dataIn1 = 32'd17
; 
32'd5897: dataIn1 = 32'd18
; 
32'd5898: dataIn1 = 32'd23
; 
32'd5899: dataIn1 = 32'd24
; 
32'd5900: dataIn1 = 32'd27
; 
32'd5901: dataIn1 = 32'd28
; 
32'd5902: dataIn1 = 32'd29
; 
32'd5903: dataIn1 = 32'd0
; 
32'd5904: dataIn1 = 32'd4
; 
32'd5905: dataIn1 = 32'd7
; 
32'd5906: dataIn1 = 32'd9
; 
32'd5907: dataIn1 = 32'd11
; 
32'd5908: dataIn1 = 32'd12
; 
32'd5909: dataIn1 = 32'd16
; 
32'd5910: dataIn1 = 32'd17
; 
32'd5911: dataIn1 = 32'd19
; 
32'd5912: dataIn1 = 32'd22
; 
32'd5913: dataIn1 = 32'd26
; 
32'd5914: dataIn1 = 32'd27
; 
32'd5915: dataIn1 = 32'd28
; 
32'd5916: dataIn1 = 32'd0
; 
32'd5917: dataIn1 = 32'd1
; 
32'd5918: dataIn1 = 32'd4
; 
32'd5919: dataIn1 = 32'd10
; 
32'd5920: dataIn1 = 32'd11
; 
32'd5921: dataIn1 = 32'd13
; 
32'd5922: dataIn1 = 32'd14
; 
32'd5923: dataIn1 = 32'd15
; 
32'd5924: dataIn1 = 32'd19
; 
32'd5925: dataIn1 = 32'd20
; 
32'd5926: dataIn1 = 32'd21
; 
32'd5927: dataIn1 = 32'd23
; 
32'd5928: dataIn1 = 32'd24
; 
32'd5929: dataIn1 = 32'd25
; 
32'd5930: dataIn1 = 32'd27
; 
32'd5931: dataIn1 = 32'd28
; 
32'd5932: dataIn1 = 32'd31
; 
32'd5933: dataIn1 = 32'd0
; 
32'd5934: dataIn1 = 32'd2
; 
32'd5935: dataIn1 = 32'd9
; 
32'd5936: dataIn1 = 32'd11
; 
32'd5937: dataIn1 = 32'd13
; 
32'd5938: dataIn1 = 32'd19
; 
32'd5939: dataIn1 = 32'd20
; 
32'd5940: dataIn1 = 32'd22
; 
32'd5941: dataIn1 = 32'd23
; 
32'd5942: dataIn1 = 32'd30
; 
32'd5943: dataIn1 = 32'd31
; 
32'd5944: dataIn1 = 32'd0
; 
32'd5945: dataIn1 = 32'd3
; 
32'd5946: dataIn1 = 32'd9
; 
32'd5947: dataIn1 = 32'd16
; 
32'd5948: dataIn1 = 32'd18
; 
32'd5949: dataIn1 = 32'd20
; 
32'd5950: dataIn1 = 32'd21
; 
32'd5951: dataIn1 = 32'd23
; 
32'd5952: dataIn1 = 32'd28
; 
32'd5953: dataIn1 = 32'd29
; 
32'd5954: dataIn1 = 32'd31
; 
32'd5955: dataIn1 = 32'd1
; 
32'd5956: dataIn1 = 32'd3
; 
32'd5957: dataIn1 = 32'd5
; 
32'd5958: dataIn1 = 32'd7
; 
32'd5959: dataIn1 = 32'd10
; 
32'd5960: dataIn1 = 32'd12
; 
32'd5961: dataIn1 = 32'd13
; 
32'd5962: dataIn1 = 32'd23
; 
32'd5963: dataIn1 = 32'd25
; 
32'd5964: dataIn1 = 32'd28
; 
32'd5965: dataIn1 = 32'd29
; 
32'd5966: dataIn1 = 32'd0
; 
32'd5967: dataIn1 = 32'd3
; 
32'd5968: dataIn1 = 32'd8
; 
32'd5969: dataIn1 = 32'd11
; 
32'd5970: dataIn1 = 32'd13
; 
32'd5971: dataIn1 = 32'd14
; 
32'd5972: dataIn1 = 32'd15
; 
32'd5973: dataIn1 = 32'd18
; 
32'd5974: dataIn1 = 32'd19
; 
32'd5975: dataIn1 = 32'd20
; 
32'd5976: dataIn1 = 32'd23
; 
32'd5977: dataIn1 = 32'd24
; 
32'd5978: dataIn1 = 32'd25
; 
32'd5979: dataIn1 = 32'd27
; 
32'd5980: dataIn1 = 32'd28
; 
32'd5981: dataIn1 = 32'd29
; 
32'd5982: dataIn1 = 32'd6
; 
32'd5983: dataIn1 = 32'd10
; 
32'd5984: dataIn1 = 32'd12
; 
32'd5985: dataIn1 = 32'd17
; 
32'd5986: dataIn1 = 32'd19
; 
32'd5987: dataIn1 = 32'd20
; 
32'd5988: dataIn1 = 32'd24
; 
32'd5989: dataIn1 = 32'd25
; 
32'd5990: dataIn1 = 32'd26
; 
32'd5991: dataIn1 = 32'd30
; 
32'd5992: dataIn1 = 32'd0
; 
32'd5993: dataIn1 = 32'd2
; 
32'd5994: dataIn1 = 32'd4
; 
32'd5995: dataIn1 = 32'd5
; 
32'd5996: dataIn1 = 32'd8
; 
32'd5997: dataIn1 = 32'd12
; 
32'd5998: dataIn1 = 32'd13
; 
32'd5999: dataIn1 = 32'd19
; 
32'd6000: dataIn1 = 32'd20
; 
32'd6001: dataIn1 = 32'd22
; 
32'd6002: dataIn1 = 32'd24
; 
32'd6003: dataIn1 = 32'd25
; 
32'd6004: dataIn1 = 32'd26
; 
32'd6005: dataIn1 = 32'd27
; 
32'd6006: dataIn1 = 32'd28
; 
32'd6007: dataIn1 = 32'd29
; 
32'd6008: dataIn1 = 32'd30
; 
32'd6009: dataIn1 = 32'd31
; 
32'd6010: dataIn1 = 32'd1
; 
32'd6011: dataIn1 = 32'd4
; 
32'd6012: dataIn1 = 32'd5
; 
32'd6013: dataIn1 = 32'd7
; 
32'd6014: dataIn1 = 32'd11
; 
32'd6015: dataIn1 = 32'd12
; 
32'd6016: dataIn1 = 32'd16
; 
32'd6017: dataIn1 = 32'd23
; 
32'd6018: dataIn1 = 32'd24
; 
32'd6019: dataIn1 = 32'd25
; 
32'd6020: dataIn1 = 32'd26
; 
32'd6021: dataIn1 = 32'd29
; 
32'd6022: dataIn1 = 32'd2
; 
32'd6023: dataIn1 = 32'd7
; 
32'd6024: dataIn1 = 32'd9
; 
32'd6025: dataIn1 = 32'd10
; 
32'd6026: dataIn1 = 32'd14
; 
32'd6027: dataIn1 = 32'd16
; 
32'd6028: dataIn1 = 32'd18
; 
32'd6029: dataIn1 = 32'd21
; 
32'd6030: dataIn1 = 32'd23
; 
32'd6031: dataIn1 = 32'd27
; 
32'd6032: dataIn1 = 32'd30
; 
32'd6033: dataIn1 = 32'd1
; 
32'd6034: dataIn1 = 32'd7
; 
32'd6035: dataIn1 = 32'd8
; 
32'd6036: dataIn1 = 32'd12
; 
32'd6037: dataIn1 = 32'd24
; 
32'd6038: dataIn1 = 32'd26
; 
32'd6039: dataIn1 = 32'd28
; 
32'd6040: dataIn1 = 32'd1
; 
32'd6041: dataIn1 = 32'd2
; 
32'd6042: dataIn1 = 32'd5
; 
32'd6043: dataIn1 = 32'd7
; 
32'd6044: dataIn1 = 32'd8
; 
32'd6045: dataIn1 = 32'd10
; 
32'd6046: dataIn1 = 32'd11
; 
32'd6047: dataIn1 = 32'd16
; 
32'd6048: dataIn1 = 32'd19
; 
32'd6049: dataIn1 = 32'd27
; 
32'd6050: dataIn1 = 32'd28
; 
32'd6051: dataIn1 = 32'd29
; 
32'd6052: dataIn1 = 32'd31
; 
32'd6053: dataIn1 = 32'd0
; 
32'd6054: dataIn1 = 32'd4
; 
32'd6055: dataIn1 = 32'd6
; 
32'd6056: dataIn1 = 32'd9
; 
32'd6057: dataIn1 = 32'd10
; 
32'd6058: dataIn1 = 32'd11
; 
32'd6059: dataIn1 = 32'd12
; 
32'd6060: dataIn1 = 32'd13
; 
32'd6061: dataIn1 = 32'd15
; 
32'd6062: dataIn1 = 32'd21
; 
32'd6063: dataIn1 = 32'd22
; 
32'd6064: dataIn1 = 32'd27
; 
32'd6065: dataIn1 = 32'd31
; 
32'd6066: dataIn1 = 32'd3
; 
32'd6067: dataIn1 = 32'd7
; 
32'd6068: dataIn1 = 32'd9
; 
32'd6069: dataIn1 = 32'd13
; 
32'd6070: dataIn1 = 32'd14
; 
32'd6071: dataIn1 = 32'd15
; 
32'd6072: dataIn1 = 32'd16
; 
32'd6073: dataIn1 = 32'd20
; 
32'd6074: dataIn1 = 32'd24
; 
32'd6075: dataIn1 = 32'd30
; 
32'd6076: dataIn1 = 32'd31
; 
32'd6077: dataIn1 = 32'd0
; 
32'd6078: dataIn1 = 32'd1
; 
32'd6079: dataIn1 = 32'd2
; 
32'd6080: dataIn1 = 32'd7
; 
32'd6081: dataIn1 = 32'd12
; 
32'd6082: dataIn1 = 32'd15
; 
32'd6083: dataIn1 = 32'd16
; 
32'd6084: dataIn1 = 32'd20
; 
32'd6085: dataIn1 = 32'd23
; 
32'd6086: dataIn1 = 32'd25
; 
32'd6087: dataIn1 = 32'd26
; 
32'd6088: dataIn1 = 32'd28
; 
32'd6089: dataIn1 = 32'd31
; 
32'd6090: dataIn1 = 32'd1
; 
32'd6091: dataIn1 = 32'd2
; 
32'd6092: dataIn1 = 32'd10
; 
32'd6093: dataIn1 = 32'd13
; 
32'd6094: dataIn1 = 32'd19
; 
32'd6095: dataIn1 = 32'd26
; 
32'd6096: dataIn1 = 32'd29
; 
32'd6097: dataIn1 = 32'd31
; 
32'd6098: dataIn1 = 32'd5
; 
32'd6099: dataIn1 = 32'd8
; 
32'd6100: dataIn1 = 32'd11
; 
32'd6101: dataIn1 = 32'd12
; 
32'd6102: dataIn1 = 32'd13
; 
32'd6103: dataIn1 = 32'd14
; 
32'd6104: dataIn1 = 32'd16
; 
32'd6105: dataIn1 = 32'd17
; 
32'd6106: dataIn1 = 32'd18
; 
32'd6107: dataIn1 = 32'd19
; 
32'd6108: dataIn1 = 32'd23
; 
32'd6109: dataIn1 = 32'd25
; 
32'd6110: dataIn1 = 32'd29
; 
32'd6111: dataIn1 = 32'd0
; 
32'd6112: dataIn1 = 32'd2
; 
32'd6113: dataIn1 = 32'd6
; 
32'd6114: dataIn1 = 32'd7
; 
32'd6115: dataIn1 = 32'd9
; 
32'd6116: dataIn1 = 32'd13
; 
32'd6117: dataIn1 = 32'd14
; 
32'd6118: dataIn1 = 32'd17
; 
32'd6119: dataIn1 = 32'd19
; 
32'd6120: dataIn1 = 32'd20
; 
32'd6121: dataIn1 = 32'd22
; 
32'd6122: dataIn1 = 32'd24
; 
32'd6123: dataIn1 = 32'd30
; 
32'd6124: dataIn1 = 32'd31
; 
32'd6125: dataIn1 = 32'd1
; 
32'd6126: dataIn1 = 32'd10
; 
32'd6127: dataIn1 = 32'd13
; 
32'd6128: dataIn1 = 32'd14
; 
32'd6129: dataIn1 = 32'd18
; 
32'd6130: dataIn1 = 32'd24
; 
32'd6131: dataIn1 = 32'd25
; 
32'd6132: dataIn1 = 32'd27
; 
32'd6133: dataIn1 = 32'd28
; 
32'd6134: dataIn1 = 32'd31
; 
32'd6135: dataIn1 = 32'd3
; 
32'd6136: dataIn1 = 32'd12
; 
32'd6137: dataIn1 = 32'd13
; 
32'd6138: dataIn1 = 32'd15
; 
32'd6139: dataIn1 = 32'd16
; 
32'd6140: dataIn1 = 32'd21
; 
32'd6141: dataIn1 = 32'd23
; 
32'd6142: dataIn1 = 32'd24
; 
32'd6143: dataIn1 = 32'd26
; 
32'd6144: dataIn1 = 32'd1
; 
32'd6145: dataIn1 = 32'd2
; 
32'd6146: dataIn1 = 32'd13
; 
32'd6147: dataIn1 = 32'd19
; 
32'd6148: dataIn1 = 32'd22
; 
32'd6149: dataIn1 = 32'd25
; 
32'd6150: dataIn1 = 32'd0
; 
32'd6151: dataIn1 = 32'd1
; 
32'd6152: dataIn1 = 32'd2
; 
32'd6153: dataIn1 = 32'd3
; 
32'd6154: dataIn1 = 32'd4
; 
32'd6155: dataIn1 = 32'd5
; 
32'd6156: dataIn1 = 32'd9
; 
32'd6157: dataIn1 = 32'd10
; 
32'd6158: dataIn1 = 32'd12
; 
32'd6159: dataIn1 = 32'd14
; 
32'd6160: dataIn1 = 32'd16
; 
32'd6161: dataIn1 = 32'd18
; 
32'd6162: dataIn1 = 32'd20
; 
32'd6163: dataIn1 = 32'd25
; 
32'd6164: dataIn1 = 32'd30
; 
32'd6165: dataIn1 = 32'd2
; 
32'd6166: dataIn1 = 32'd4
; 
32'd6167: dataIn1 = 32'd5
; 
32'd6168: dataIn1 = 32'd7
; 
32'd6169: dataIn1 = 32'd11
; 
32'd6170: dataIn1 = 32'd12
; 
32'd6171: dataIn1 = 32'd14
; 
32'd6172: dataIn1 = 32'd15
; 
32'd6173: dataIn1 = 32'd16
; 
32'd6174: dataIn1 = 32'd17
; 
32'd6175: dataIn1 = 32'd20
; 
32'd6176: dataIn1 = 32'd26
; 
32'd6177: dataIn1 = 32'd29
; 
32'd6178: dataIn1 = 32'd30
; 
32'd6179: dataIn1 = 32'd1
; 
32'd6180: dataIn1 = 32'd4
; 
32'd6181: dataIn1 = 32'd5
; 
32'd6182: dataIn1 = 32'd6
; 
32'd6183: dataIn1 = 32'd7
; 
32'd6184: dataIn1 = 32'd14
; 
32'd6185: dataIn1 = 32'd15
; 
32'd6186: dataIn1 = 32'd16
; 
32'd6187: dataIn1 = 32'd20
; 
32'd6188: dataIn1 = 32'd22
; 
32'd6189: dataIn1 = 32'd24
; 
32'd6190: dataIn1 = 32'd25
; 
32'd6191: dataIn1 = 32'd28
; 
32'd6192: dataIn1 = 32'd29
; 
32'd6193: dataIn1 = 32'd0
; 
32'd6194: dataIn1 = 32'd4
; 
32'd6195: dataIn1 = 32'd5
; 
32'd6196: dataIn1 = 32'd8
; 
32'd6197: dataIn1 = 32'd11
; 
32'd6198: dataIn1 = 32'd12
; 
32'd6199: dataIn1 = 32'd16
; 
32'd6200: dataIn1 = 32'd18
; 
32'd6201: dataIn1 = 32'd20
; 
32'd6202: dataIn1 = 32'd21
; 
32'd6203: dataIn1 = 32'd26
; 
32'd6204: dataIn1 = 32'd27
; 
32'd6205: dataIn1 = 32'd28
; 
32'd6206: dataIn1 = 32'd29
; 
32'd6207: dataIn1 = 32'd30
; 
32'd6208: dataIn1 = 32'd0
; 
32'd6209: dataIn1 = 32'd1
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd90; 
32'd3: dataIn2 = 32'd51; 
32'd4: dataIn2 = 32'd93; 
32'd5: dataIn2 = 32'd89; 
32'd6: dataIn2 = 32'd62; 
32'd7: dataIn2 = 32'd6; 
32'd8: dataIn2 = 32'd50; 
32'd9: dataIn2 = 32'd21; 
32'd10: dataIn2 = 32'd96; 
32'd11: dataIn2 = 32'd33; 
32'd12: dataIn2 = 32'd49; 
32'd13: dataIn2 = 32'd61; 
32'd14: dataIn2 = 32'd90; 
32'd15: dataIn2 = 32'd33; 
32'd16: dataIn2 = 32'd81; 
32'd17: dataIn2 = 32'd44; 
32'd18: dataIn2 = 32'd55; 
32'd19: dataIn2 = 32'd61; 
32'd20: dataIn2 = 32'd54; 
32'd21: dataIn2 = 32'd34; 
32'd22: dataIn2 = 32'd60; 
32'd23: dataIn2 = 32'd5; 
32'd24: dataIn2 = 32'd100; 
32'd25: dataIn2 = 32'd23; 
32'd26: dataIn2 = 32'd81; 
32'd27: dataIn2 = 32'd97; 
32'd28: dataIn2 = 32'd23; 
32'd29: dataIn2 = 32'd73; 
32'd30: dataIn2 = 32'd48; 
32'd31: dataIn2 = 32'd36; 
32'd32: dataIn2 = 32'd15; 
32'd33: dataIn2 = 32'd8; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd170: dataIn2 = 32'd59; 
32'd171: dataIn2 = 32'd66; 
32'd172: dataIn2 = 32'd50; 
32'd173: dataIn2 = 32'd31; 
32'd174: dataIn2 = 32'd34; 
32'd175: dataIn2 = 32'd98; 
32'd176: dataIn2 = 32'd51; 
32'd177: dataIn2 = 32'd35; 
32'd178: dataIn2 = 32'd18; 
32'd179: dataIn2 = 32'd21; 
32'd180: dataIn2 = 32'd66; 
32'd181: dataIn2 = 32'd63; 
32'd182: dataIn2 = 32'd91; 
32'd183: dataIn2 = 32'd98; 
32'd184: dataIn2 = 32'd24; 
32'd185: dataIn2 = 32'd58; 
32'd186: dataIn2 = 32'd80; 
32'd187: dataIn2 = 32'd47; 
32'd188: dataIn2 = 32'd77; 
32'd189: dataIn2 = 32'd57; 
32'd190: dataIn2 = 32'd95; 
32'd191: dataIn2 = 32'd5; 
32'd192: dataIn2 = 32'd39; 
32'd193: dataIn2 = 32'd87; 
32'd194: dataIn2 = 32'd25; 
32'd195: dataIn2 = 32'd78; 
32'd196: dataIn2 = 32'd61; 
32'd197: dataIn2 = 32'd90; 
32'd198: dataIn2 = 32'd85; 
32'd199: dataIn2 = 32'd29; 
32'd200: dataIn2 = 32'd1; 
32'd201: dataIn2 = 32'd5; 
32'd202: dataIn2 = 32'd99; 
32'd203: dataIn2 = 32'd95; 
32'd204: dataIn2 = 32'd98; 
32'd205: dataIn2 = 32'd39; 
32'd206: dataIn2 = 32'd14; 
32'd207: dataIn2 = 32'd25; 
32'd208: dataIn2 = 32'd85; 
32'd209: dataIn2 = 32'd50; 
32'd210: dataIn2 = 32'd67; 
32'd211: dataIn2 = 32'd55; 
32'd212: dataIn2 = 32'd73; 
32'd213: dataIn2 = 32'd12; 
32'd214: dataIn2 = 32'd75; 
32'd215: dataIn2 = 32'd51; 
32'd216: dataIn2 = 32'd76; 
32'd217: dataIn2 = 32'd73; 
32'd218: dataIn2 = 32'd4; 
32'd219: dataIn2 = 32'd1; 
32'd220: dataIn2 = 32'd56; 
32'd221: dataIn2 = 32'd69; 
32'd222: dataIn2 = 32'd14; 
32'd223: dataIn2 = 32'd40; 
32'd224: dataIn2 = 32'd49; 
32'd225: dataIn2 = 32'd72; 
32'd226: dataIn2 = 32'd85; 
32'd227: dataIn2 = 32'd58; 
32'd228: dataIn2 = 32'd29; 
32'd229: dataIn2 = 32'd48; 
32'd230: dataIn2 = 32'd52; 
32'd231: dataIn2 = 32'd78; 
32'd232: dataIn2 = 32'd34; 
32'd233: dataIn2 = 32'd80; 
32'd234: dataIn2 = 32'd56; 
32'd235: dataIn2 = 32'd19; 
32'd236: dataIn2 = 32'd97; 
32'd237: dataIn2 = 32'd48; 
32'd238: dataIn2 = 32'd43; 
32'd239: dataIn2 = 32'd13; 
32'd240: dataIn2 = 32'd93; 
32'd241: dataIn2 = 32'd52; 
32'd242: dataIn2 = 32'd13; 
32'd243: dataIn2 = 32'd11; 
32'd244: dataIn2 = 32'd95; 
32'd245: dataIn2 = 32'd52; 
32'd246: dataIn2 = 32'd75; 
32'd247: dataIn2 = 32'd35; 
32'd248: dataIn2 = 32'd20; 
32'd249: dataIn2 = 32'd35; 
32'd250: dataIn2 = 32'd94; 
32'd251: dataIn2 = 32'd53; 
32'd252: dataIn2 = 32'd7; 
32'd253: dataIn2 = 32'd74; 
32'd254: dataIn2 = 32'd3; 
32'd255: dataIn2 = 32'd47; 
32'd256: dataIn2 = 32'd79; 
32'd257: dataIn2 = 32'd64; 
32'd258: dataIn2 = 32'd59; 
32'd259: dataIn2 = 32'd33; 
32'd260: dataIn2 = 32'd3; 
32'd261: dataIn2 = 32'd32; 
32'd262: dataIn2 = 32'd15; 
32'd263: dataIn2 = 32'd73; 
32'd264: dataIn2 = 32'd27; 
32'd265: dataIn2 = 32'd12; 
32'd266: dataIn2 = 32'd72; 
32'd267: dataIn2 = 32'd76; 
32'd268: dataIn2 = 32'd74; 
32'd269: dataIn2 = 32'd54; 
32'd270: dataIn2 = 32'd30; 
32'd271: dataIn2 = 32'd40; 
32'd272: dataIn2 = 32'd62; 
32'd273: dataIn2 = 32'd20; 
32'd274: dataIn2 = 32'd85; 
32'd275: dataIn2 = 32'd36; 
32'd276: dataIn2 = 32'd96; 
32'd277: dataIn2 = 32'd35; 
32'd278: dataIn2 = 32'd91; 
32'd279: dataIn2 = 32'd35; 
32'd280: dataIn2 = 32'd17; 
32'd281: dataIn2 = 32'd18; 
32'd282: dataIn2 = 32'd24; 
32'd283: dataIn2 = 32'd13; 
32'd284: dataIn2 = 32'd86; 
32'd285: dataIn2 = 32'd26; 
32'd286: dataIn2 = 32'd1; 
32'd287: dataIn2 = 32'd41; 
32'd288: dataIn2 = 32'd39; 
32'd289: dataIn2 = 32'd7; 
32'd290: dataIn2 = 32'd34; 
32'd291: dataIn2 = 32'd22; 
32'd292: dataIn2 = 32'd49; 
32'd293: dataIn2 = 32'd96; 
32'd294: dataIn2 = 32'd19; 
32'd295: dataIn2 = 32'd51; 
32'd296: dataIn2 = 32'd64; 
32'd297: dataIn2 = 32'd99; 
32'd298: dataIn2 = 32'd54; 
32'd299: dataIn2 = 32'd54; 
32'd300: dataIn2 = 32'd67; 
32'd301: dataIn2 = 32'd37; 
32'd302: dataIn2 = 32'd51; 
32'd303: dataIn2 = 32'd1; 
32'd304: dataIn2 = 32'd21; 
32'd305: dataIn2 = 32'd88; 
32'd306: dataIn2 = 32'd80; 
32'd307: dataIn2 = 32'd47; 
32'd308: dataIn2 = 32'd49; 
32'd309: dataIn2 = 32'd35; 
32'd310: dataIn2 = 32'd4; 
32'd311: dataIn2 = 32'd45; 
32'd312: dataIn2 = 32'd7; 
32'd313: dataIn2 = 32'd42; 
32'd314: dataIn2 = 32'd17; 
32'd315: dataIn2 = 32'd89; 
32'd316: dataIn2 = 32'd0; 
32'd317: dataIn2 = 32'd63; 
32'd318: dataIn2 = 32'd92; 
32'd319: dataIn2 = 32'd41; 
32'd320: dataIn2 = 32'd49; 
32'd321: dataIn2 = 32'd29; 
32'd322: dataIn2 = 32'd69; 
32'd323: dataIn2 = 32'd74; 
32'd324: dataIn2 = 32'd59; 
32'd325: dataIn2 = 32'd72; 
32'd326: dataIn2 = 32'd89; 
32'd327: dataIn2 = 32'd15; 
32'd328: dataIn2 = 32'd42; 
32'd329: dataIn2 = 32'd76; 
32'd330: dataIn2 = 32'd4; 
32'd331: dataIn2 = 32'd63; 
32'd332: dataIn2 = 32'd58; 
32'd333: dataIn2 = 32'd61; 
32'd334: dataIn2 = 32'd22; 
32'd335: dataIn2 = 32'd13; 
32'd336: dataIn2 = 32'd57; 
32'd337: dataIn2 = 32'd97; 
32'd338: dataIn2 = 32'd91; 
32'd339: dataIn2 = 32'd33; 
32'd340: dataIn2 = 32'd66; 
32'd341: dataIn2 = 32'd10; 
32'd342: dataIn2 = 32'd24; 
32'd343: dataIn2 = 32'd43; 
32'd344: dataIn2 = 32'd89; 
32'd345: dataIn2 = 32'd65; 
32'd346: dataIn2 = 32'd97; 
32'd347: dataIn2 = 32'd96; 
32'd348: dataIn2 = 32'd71; 
32'd349: dataIn2 = 32'd93; 
32'd350: dataIn2 = 32'd17; 
32'd351: dataIn2 = 32'd26; 
32'd352: dataIn2 = 32'd34; 
32'd353: dataIn2 = 32'd95; 
32'd354: dataIn2 = 32'd25; 
32'd355: dataIn2 = 32'd33; 
32'd356: dataIn2 = 32'd45; 
32'd357: dataIn2 = 32'd25; 
32'd358: dataIn2 = 32'd72; 
32'd359: dataIn2 = 32'd90; 
32'd360: dataIn2 = 32'd31; 
32'd361: dataIn2 = 32'd33; 
32'd362: dataIn2 = 32'd33; 
32'd363: dataIn2 = 32'd49; 
32'd364: dataIn2 = 32'd72; 
32'd365: dataIn2 = 32'd16; 
32'd366: dataIn2 = 32'd22; 
32'd367: dataIn2 = 32'd35; 
32'd368: dataIn2 = 32'd77; 
32'd369: dataIn2 = 32'd44; 
32'd370: dataIn2 = 32'd36; 
32'd371: dataIn2 = 32'd86; 
32'd372: dataIn2 = 32'd98; 
32'd373: dataIn2 = 32'd4; 
32'd374: dataIn2 = 32'd87; 
32'd375: dataIn2 = 32'd84; 
32'd376: dataIn2 = 32'd30; 
32'd377: dataIn2 = 32'd51; 
32'd378: dataIn2 = 32'd79; 
32'd379: dataIn2 = 32'd44; 
32'd380: dataIn2 = 32'd83; 
32'd381: dataIn2 = 32'd35; 
32'd382: dataIn2 = 32'd5; 
32'd383: dataIn2 = 32'd38; 
32'd384: dataIn2 = 32'd87; 
32'd385: dataIn2 = 32'd93; 
32'd386: dataIn2 = 32'd28; 
32'd387: dataIn2 = 32'd100; 
32'd388: dataIn2 = 32'd20; 
32'd389: dataIn2 = 32'd16; 
32'd390: dataIn2 = 32'd44; 
32'd391: dataIn2 = 32'd75; 
32'd392: dataIn2 = 32'd41; 
32'd393: dataIn2 = 32'd11; 
32'd394: dataIn2 = 32'd24; 
32'd395: dataIn2 = 32'd98; 
32'd396: dataIn2 = 32'd23; 
32'd397: dataIn2 = 32'd30; 
32'd398: dataIn2 = 32'd30; 
32'd399: dataIn2 = 32'd67; 
32'd400: dataIn2 = 32'd49; 
32'd401: dataIn2 = 32'd65; 
32'd402: dataIn2 = 32'd38; 
32'd403: dataIn2 = 32'd41; 
32'd404: dataIn2 = 32'd20; 
32'd405: dataIn2 = 32'd10; 
32'd406: dataIn2 = 32'd14; 
32'd407: dataIn2 = 32'd80; 
32'd408: dataIn2 = 32'd3; 
32'd409: dataIn2 = 32'd62; 
32'd410: dataIn2 = 32'd58; 
32'd411: dataIn2 = 32'd91; 
32'd412: dataIn2 = 32'd11; 
32'd413: dataIn2 = 32'd83; 
32'd414: dataIn2 = 32'd1; 
32'd415: dataIn2 = 32'd36; 
32'd416: dataIn2 = 32'd46; 
32'd417: dataIn2 = 32'd17; 
32'd418: dataIn2 = 32'd25; 
32'd419: dataIn2 = 32'd51; 
32'd420: dataIn2 = 32'd17; 
32'd421: dataIn2 = 32'd94; 
32'd422: dataIn2 = 32'd35; 
32'd423: dataIn2 = 32'd100; 
32'd424: dataIn2 = 32'd41; 
32'd425: dataIn2 = 32'd3; 
32'd426: dataIn2 = 32'd44; 
32'd427: dataIn2 = 32'd45; 
32'd428: dataIn2 = 32'd17; 
32'd429: dataIn2 = 32'd42; 
32'd430: dataIn2 = 32'd89; 
32'd431: dataIn2 = 32'd1; 
32'd432: dataIn2 = 32'd35; 
32'd433: dataIn2 = 32'd90; 
32'd434: dataIn2 = 32'd7; 
32'd435: dataIn2 = 32'd98; 
32'd436: dataIn2 = 32'd12; 
32'd437: dataIn2 = 32'd36; 
32'd438: dataIn2 = 32'd40; 
32'd439: dataIn2 = 32'd79; 
32'd440: dataIn2 = 32'd33; 
32'd441: dataIn2 = 32'd30; 
32'd442: dataIn2 = 32'd25; 
32'd443: dataIn2 = 32'd91; 
32'd444: dataIn2 = 32'd64; 
32'd445: dataIn2 = 32'd65; 
32'd446: dataIn2 = 32'd98; 
32'd447: dataIn2 = 32'd15; 
32'd448: dataIn2 = 32'd15; 
32'd449: dataIn2 = 32'd71; 
32'd450: dataIn2 = 32'd25; 
32'd451: dataIn2 = 32'd34; 
32'd452: dataIn2 = 32'd97; 
32'd453: dataIn2 = 32'd5; 
32'd454: dataIn2 = 32'd84; 
32'd455: dataIn2 = 32'd51; 
32'd456: dataIn2 = 32'd65; 
32'd457: dataIn2 = 32'd51; 
32'd458: dataIn2 = 32'd29; 
32'd459: dataIn2 = 32'd58; 
32'd460: dataIn2 = 32'd89; 
32'd461: dataIn2 = 32'd37; 
32'd462: dataIn2 = 32'd52; 
32'd463: dataIn2 = 32'd100; 
32'd464: dataIn2 = 32'd79; 
32'd465: dataIn2 = 32'd77; 
32'd466: dataIn2 = 32'd94; 
32'd467: dataIn2 = 32'd95; 
32'd468: dataIn2 = 32'd28; 
32'd469: dataIn2 = 32'd81; 
32'd470: dataIn2 = 32'd72; 
32'd471: dataIn2 = 32'd9; 
32'd472: dataIn2 = 32'd38; 
32'd473: dataIn2 = 32'd60; 
32'd474: dataIn2 = 32'd75; 
32'd475: dataIn2 = 32'd94; 
32'd476: dataIn2 = 32'd63; 
32'd477: dataIn2 = 32'd2; 
32'd478: dataIn2 = 32'd88; 
32'd479: dataIn2 = 32'd81; 
32'd480: dataIn2 = 32'd96; 
32'd481: dataIn2 = 32'd20; 
32'd482: dataIn2 = 32'd74; 
32'd483: dataIn2 = 32'd93; 
32'd484: dataIn2 = 32'd39; 
32'd485: dataIn2 = 32'd18; 
32'd486: dataIn2 = 32'd70; 
32'd487: dataIn2 = 32'd79; 
32'd488: dataIn2 = 32'd68; 
32'd489: dataIn2 = 32'd98; 
32'd490: dataIn2 = 32'd24; 
32'd491: dataIn2 = 32'd70; 
32'd492: dataIn2 = 32'd13; 
32'd493: dataIn2 = 32'd5; 
32'd494: dataIn2 = 32'd85; 
32'd495: dataIn2 = 32'd43; 
32'd496: dataIn2 = 32'd42; 
32'd497: dataIn2 = 32'd39; 
32'd498: dataIn2 = 32'd11; 
32'd499: dataIn2 = 32'd95; 
32'd500: dataIn2 = 32'd100; 
32'd501: dataIn2 = 32'd99; 
32'd502: dataIn2 = 32'd32; 
32'd503: dataIn2 = 32'd24; 
32'd504: dataIn2 = 32'd36; 
32'd505: dataIn2 = 32'd0; 
32'd506: dataIn2 = 32'd67; 
32'd507: dataIn2 = 32'd75; 
32'd508: dataIn2 = 32'd93; 
32'd509: dataIn2 = 32'd7; 
32'd510: dataIn2 = 32'd39; 
32'd511: dataIn2 = 32'd22; 
32'd512: dataIn2 = 32'd34; 
32'd513: dataIn2 = 32'd90; 
32'd514: dataIn2 = 32'd50; 
32'd515: dataIn2 = 32'd90; 
32'd516: dataIn2 = 32'd73; 
32'd517: dataIn2 = 32'd60; 
32'd518: dataIn2 = 32'd89; 
32'd519: dataIn2 = 32'd69; 
32'd520: dataIn2 = 32'd29; 
32'd521: dataIn2 = 32'd48; 
32'd522: dataIn2 = 32'd11; 
32'd523: dataIn2 = 32'd78; 
32'd524: dataIn2 = 32'd71; 
32'd525: dataIn2 = 32'd74; 
32'd526: dataIn2 = 32'd63; 
32'd527: dataIn2 = 32'd70; 
32'd528: dataIn2 = 32'd15; 
32'd529: dataIn2 = 32'd36; 
32'd530: dataIn2 = 32'd27; 
32'd531: dataIn2 = 32'd42; 
32'd532: dataIn2 = 32'd30; 
32'd533: dataIn2 = 32'd9; 
32'd534: dataIn2 = 32'd34; 
32'd535: dataIn2 = 32'd13; 
32'd536: dataIn2 = 32'd42; 
32'd537: dataIn2 = 32'd37; 
32'd538: dataIn2 = 32'd51; 
32'd539: dataIn2 = 32'd63; 
32'd540: dataIn2 = 32'd19; 
32'd541: dataIn2 = 32'd12; 
32'd542: dataIn2 = 32'd71; 
32'd543: dataIn2 = 32'd90; 
32'd544: dataIn2 = 32'd28; 
32'd545: dataIn2 = 32'd26; 
32'd546: dataIn2 = 32'd95; 
32'd547: dataIn2 = 32'd25; 
32'd548: dataIn2 = 32'd38; 
32'd549: dataIn2 = 32'd89; 
32'd550: dataIn2 = 32'd3; 
32'd551: dataIn2 = 32'd27; 
32'd552: dataIn2 = 32'd41; 
32'd553: dataIn2 = 32'd60; 
32'd554: dataIn2 = 32'd36; 
32'd555: dataIn2 = 32'd95; 
32'd556: dataIn2 = 32'd60; 
32'd557: dataIn2 = 32'd88; 
32'd558: dataIn2 = 32'd17; 
32'd559: dataIn2 = 32'd72; 
32'd560: dataIn2 = 32'd92; 
32'd561: dataIn2 = 32'd43; 
32'd562: dataIn2 = 32'd19; 
32'd563: dataIn2 = 32'd19; 
32'd564: dataIn2 = 32'd16; 
32'd565: dataIn2 = 32'd37; 
32'd566: dataIn2 = 32'd2; 
32'd567: dataIn2 = 32'd53; 
32'd568: dataIn2 = 32'd80; 
32'd569: dataIn2 = 32'd90; 
32'd570: dataIn2 = 32'd45; 
32'd571: dataIn2 = 32'd42; 
32'd572: dataIn2 = 32'd3; 
32'd573: dataIn2 = 32'd94; 
32'd574: dataIn2 = 32'd3; 
32'd575: dataIn2 = 32'd27; 
32'd576: dataIn2 = 32'd25; 
32'd577: dataIn2 = 32'd62; 
32'd578: dataIn2 = 32'd59; 
32'd579: dataIn2 = 32'd73; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_32_60.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
