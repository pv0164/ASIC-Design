//64x64 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 2867 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd330 ; 
  wdata_col_base = 32'd31970 ; 
  row_base = 32'd348370 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #302000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd348370: dataIn1 = 32'd0
; 
32'd348371: dataIn1 = 32'd43
; 
32'd348372: dataIn1 = 32'd84
; 
32'd348373: dataIn1 = 32'd127
; 
32'd348374: dataIn1 = 32'd167
; 
32'd348375: dataIn1 = 32'd213
; 
32'd348376: dataIn1 = 32'd258
; 
32'd348377: dataIn1 = 32'd301
; 
32'd348378: dataIn1 = 32'd350
; 
32'd348379: dataIn1 = 32'd385
; 
32'd348380: dataIn1 = 32'd432
; 
32'd348381: dataIn1 = 32'd482
; 
32'd348382: dataIn1 = 32'd524
; 
32'd348383: dataIn1 = 32'd565
; 
32'd348384: dataIn1 = 32'd605
; 
32'd348385: dataIn1 = 32'd650
; 
32'd348386: dataIn1 = 32'd691
; 
32'd348387: dataIn1 = 32'd742
; 
32'd348388: dataIn1 = 32'd782
; 
32'd348389: dataIn1 = 32'd826
; 
32'd348390: dataIn1 = 32'd874
; 
32'd348391: dataIn1 = 32'd916
; 
32'd348392: dataIn1 = 32'd964
; 
32'd348393: dataIn1 = 32'd1007
; 
32'd348394: dataIn1 = 32'd1054
; 
32'd348395: dataIn1 = 32'd1102
; 
32'd348396: dataIn1 = 32'd1145
; 
32'd348397: dataIn1 = 32'd1193
; 
32'd348398: dataIn1 = 32'd1234
; 
32'd348399: dataIn1 = 32'd1282
; 
32'd348400: dataIn1 = 32'd1327
; 
32'd348401: dataIn1 = 32'd1371
; 
32'd348402: dataIn1 = 32'd1413
; 
32'd348403: dataIn1 = 32'd1448
; 
32'd348404: dataIn1 = 32'd1492
; 
32'd348405: dataIn1 = 32'd1534
; 
32'd348406: dataIn1 = 32'd1578
; 
32'd348407: dataIn1 = 32'd1624
; 
32'd348408: dataIn1 = 32'd1668
; 
32'd348409: dataIn1 = 32'd1709
; 
32'd348410: dataIn1 = 32'd1753
; 
32'd348411: dataIn1 = 32'd1797
; 
32'd348412: dataIn1 = 32'd1841
; 
32'd348413: dataIn1 = 32'd1885
; 
32'd348414: dataIn1 = 32'd1927
; 
32'd348415: dataIn1 = 32'd1964
; 
32'd348416: dataIn1 = 32'd2010
; 
32'd348417: dataIn1 = 32'd2053
; 
32'd348418: dataIn1 = 32'd2098
; 
32'd348419: dataIn1 = 32'd2140
; 
32'd348420: dataIn1 = 32'd2182
; 
32'd348421: dataIn1 = 32'd2222
; 
32'd348422: dataIn1 = 32'd2264
; 
32'd348423: dataIn1 = 32'd2306
; 
32'd348424: dataIn1 = 32'd2350
; 
32'd348425: dataIn1 = 32'd2393
; 
32'd348426: dataIn1 = 32'd2434
; 
32'd348427: dataIn1 = 32'd2485
; 
32'd348428: dataIn1 = 32'd2522
; 
32'd348429: dataIn1 = 32'd2562
; 
32'd348430: dataIn1 = 32'd2609
; 
32'd348431: dataIn1 = 32'd2650
; 
32'd348432: dataIn1 = 32'd2692
; 
32'd348433: dataIn1 = 32'd2736
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd31970: dataIn1 = 32'd0
; 
32'd31971: dataIn1 = 32'd43
; 
32'd31972: dataIn1 = 32'd84
; 
32'd31973: dataIn1 = 32'd127
; 
32'd31974: dataIn1 = 32'd167
; 
32'd31975: dataIn1 = 32'd213
; 
32'd31976: dataIn1 = 32'd258
; 
32'd31977: dataIn1 = 32'd301
; 
32'd31978: dataIn1 = 32'd350
; 
32'd31979: dataIn1 = 32'd385
; 
32'd31980: dataIn1 = 32'd432
; 
32'd31981: dataIn1 = 32'd482
; 
32'd31982: dataIn1 = 32'd524
; 
32'd31983: dataIn1 = 32'd565
; 
32'd31984: dataIn1 = 32'd605
; 
32'd31985: dataIn1 = 32'd650
; 
32'd31986: dataIn1 = 32'd691
; 
32'd31987: dataIn1 = 32'd742
; 
32'd31988: dataIn1 = 32'd782
; 
32'd31989: dataIn1 = 32'd826
; 
32'd31990: dataIn1 = 32'd874
; 
32'd31991: dataIn1 = 32'd916
; 
32'd31992: dataIn1 = 32'd964
; 
32'd31993: dataIn1 = 32'd1007
; 
32'd31994: dataIn1 = 32'd1054
; 
32'd31995: dataIn1 = 32'd1102
; 
32'd31996: dataIn1 = 32'd1145
; 
32'd31997: dataIn1 = 32'd1193
; 
32'd31998: dataIn1 = 32'd1234
; 
32'd31999: dataIn1 = 32'd1282
; 
32'd32000: dataIn1 = 32'd1327
; 
32'd32001: dataIn1 = 32'd1371
; 
32'd32002: dataIn1 = 32'd1413
; 
32'd32003: dataIn1 = 32'd1448
; 
32'd32004: dataIn1 = 32'd1492
; 
32'd32005: dataIn1 = 32'd1534
; 
32'd32006: dataIn1 = 32'd1578
; 
32'd32007: dataIn1 = 32'd1624
; 
32'd32008: dataIn1 = 32'd1668
; 
32'd32009: dataIn1 = 32'd1709
; 
32'd32010: dataIn1 = 32'd1753
; 
32'd32011: dataIn1 = 32'd1797
; 
32'd32012: dataIn1 = 32'd1841
; 
32'd32013: dataIn1 = 32'd1885
; 
32'd32014: dataIn1 = 32'd1927
; 
32'd32015: dataIn1 = 32'd1964
; 
32'd32016: dataIn1 = 32'd2010
; 
32'd32017: dataIn1 = 32'd2053
; 
32'd32018: dataIn1 = 32'd2098
; 
32'd32019: dataIn1 = 32'd2140
; 
32'd32020: dataIn1 = 32'd2182
; 
32'd32021: dataIn1 = 32'd2222
; 
32'd32022: dataIn1 = 32'd2264
; 
32'd32023: dataIn1 = 32'd2306
; 
32'd32024: dataIn1 = 32'd2350
; 
32'd32025: dataIn1 = 32'd2393
; 
32'd32026: dataIn1 = 32'd2434
; 
32'd32027: dataIn1 = 32'd2485
; 
32'd32028: dataIn1 = 32'd2522
; 
32'd32029: dataIn1 = 32'd2562
; 
32'd32030: dataIn1 = 32'd2609
; 
32'd32031: dataIn1 = 32'd2650
; 
32'd32032: dataIn1 = 32'd2692
; 
32'd32033: dataIn1 = 32'd2736
; 
32'd32034: dataIn1 = 32'd2773
; 
32'd32035: dataIn1 = 32'd0
; 
32'd32036: dataIn1 = 32'd1
; 
32'd32037: dataIn1 = 32'd3
; 
32'd32038: dataIn1 = 32'd4
; 
32'd32039: dataIn1 = 32'd5
; 
32'd32040: dataIn1 = 32'd6
; 
32'd32041: dataIn1 = 32'd7
; 
32'd32042: dataIn1 = 32'd8
; 
32'd32043: dataIn1 = 32'd9
; 
32'd32044: dataIn1 = 32'd10
; 
32'd32045: dataIn1 = 32'd11
; 
32'd32046: dataIn1 = 32'd13
; 
32'd32047: dataIn1 = 32'd14
; 
32'd32048: dataIn1 = 32'd16
; 
32'd32049: dataIn1 = 32'd17
; 
32'd32050: dataIn1 = 32'd18
; 
32'd32051: dataIn1 = 32'd19
; 
32'd32052: dataIn1 = 32'd20
; 
32'd32053: dataIn1 = 32'd21
; 
32'd32054: dataIn1 = 32'd22
; 
32'd32055: dataIn1 = 32'd23
; 
32'd32056: dataIn1 = 32'd26
; 
32'd32057: dataIn1 = 32'd27
; 
32'd32058: dataIn1 = 32'd28
; 
32'd32059: dataIn1 = 32'd29
; 
32'd32060: dataIn1 = 32'd33
; 
32'd32061: dataIn1 = 32'd34
; 
32'd32062: dataIn1 = 32'd39
; 
32'd32063: dataIn1 = 32'd40
; 
32'd32064: dataIn1 = 32'd42
; 
32'd32065: dataIn1 = 32'd44
; 
32'd32066: dataIn1 = 32'd45
; 
32'd32067: dataIn1 = 32'd47
; 
32'd32068: dataIn1 = 32'd48
; 
32'd32069: dataIn1 = 32'd49
; 
32'd32070: dataIn1 = 32'd51
; 
32'd32071: dataIn1 = 32'd52
; 
32'd32072: dataIn1 = 32'd53
; 
32'd32073: dataIn1 = 32'd54
; 
32'd32074: dataIn1 = 32'd56
; 
32'd32075: dataIn1 = 32'd57
; 
32'd32076: dataIn1 = 32'd61
; 
32'd32077: dataIn1 = 32'd63
; 
32'd32078: dataIn1 = 32'd1
; 
32'd32079: dataIn1 = 32'd2
; 
32'd32080: dataIn1 = 32'd3
; 
32'd32081: dataIn1 = 32'd5
; 
32'd32082: dataIn1 = 32'd7
; 
32'd32083: dataIn1 = 32'd8
; 
32'd32084: dataIn1 = 32'd9
; 
32'd32085: dataIn1 = 32'd10
; 
32'd32086: dataIn1 = 32'd11
; 
32'd32087: dataIn1 = 32'd13
; 
32'd32088: dataIn1 = 32'd14
; 
32'd32089: dataIn1 = 32'd15
; 
32'd32090: dataIn1 = 32'd18
; 
32'd32091: dataIn1 = 32'd23
; 
32'd32092: dataIn1 = 32'd24
; 
32'd32093: dataIn1 = 32'd25
; 
32'd32094: dataIn1 = 32'd26
; 
32'd32095: dataIn1 = 32'd30
; 
32'd32096: dataIn1 = 32'd31
; 
32'd32097: dataIn1 = 32'd32
; 
32'd32098: dataIn1 = 32'd33
; 
32'd32099: dataIn1 = 32'd35
; 
32'd32100: dataIn1 = 32'd36
; 
32'd32101: dataIn1 = 32'd37
; 
32'd32102: dataIn1 = 32'd38
; 
32'd32103: dataIn1 = 32'd41
; 
32'd32104: dataIn1 = 32'd42
; 
32'd32105: dataIn1 = 32'd43
; 
32'd32106: dataIn1 = 32'd44
; 
32'd32107: dataIn1 = 32'd45
; 
32'd32108: dataIn1 = 32'd46
; 
32'd32109: dataIn1 = 32'd47
; 
32'd32110: dataIn1 = 32'd48
; 
32'd32111: dataIn1 = 32'd49
; 
32'd32112: dataIn1 = 32'd50
; 
32'd32113: dataIn1 = 32'd51
; 
32'd32114: dataIn1 = 32'd53
; 
32'd32115: dataIn1 = 32'd57
; 
32'd32116: dataIn1 = 32'd58
; 
32'd32117: dataIn1 = 32'd59
; 
32'd32118: dataIn1 = 32'd63
; 
32'd32119: dataIn1 = 32'd0
; 
32'd32120: dataIn1 = 32'd1
; 
32'd32121: dataIn1 = 32'd2
; 
32'd32122: dataIn1 = 32'd4
; 
32'd32123: dataIn1 = 32'd5
; 
32'd32124: dataIn1 = 32'd6
; 
32'd32125: dataIn1 = 32'd8
; 
32'd32126: dataIn1 = 32'd10
; 
32'd32127: dataIn1 = 32'd11
; 
32'd32128: dataIn1 = 32'd13
; 
32'd32129: dataIn1 = 32'd14
; 
32'd32130: dataIn1 = 32'd15
; 
32'd32131: dataIn1 = 32'd16
; 
32'd32132: dataIn1 = 32'd19
; 
32'd32133: dataIn1 = 32'd20
; 
32'd32134: dataIn1 = 32'd21
; 
32'd32135: dataIn1 = 32'd22
; 
32'd32136: dataIn1 = 32'd23
; 
32'd32137: dataIn1 = 32'd26
; 
32'd32138: dataIn1 = 32'd27
; 
32'd32139: dataIn1 = 32'd29
; 
32'd32140: dataIn1 = 32'd31
; 
32'd32141: dataIn1 = 32'd33
; 
32'd32142: dataIn1 = 32'd35
; 
32'd32143: dataIn1 = 32'd37
; 
32'd32144: dataIn1 = 32'd38
; 
32'd32145: dataIn1 = 32'd39
; 
32'd32146: dataIn1 = 32'd40
; 
32'd32147: dataIn1 = 32'd41
; 
32'd32148: dataIn1 = 32'd43
; 
32'd32149: dataIn1 = 32'd44
; 
32'd32150: dataIn1 = 32'd45
; 
32'd32151: dataIn1 = 32'd46
; 
32'd32152: dataIn1 = 32'd48
; 
32'd32153: dataIn1 = 32'd49
; 
32'd32154: dataIn1 = 32'd50
; 
32'd32155: dataIn1 = 32'd51
; 
32'd32156: dataIn1 = 32'd53
; 
32'd32157: dataIn1 = 32'd55
; 
32'd32158: dataIn1 = 32'd58
; 
32'd32159: dataIn1 = 32'd60
; 
32'd32160: dataIn1 = 32'd61
; 
32'd32161: dataIn1 = 32'd63
; 
32'd32162: dataIn1 = 32'd1
; 
32'd32163: dataIn1 = 32'd3
; 
32'd32164: dataIn1 = 32'd4
; 
32'd32165: dataIn1 = 32'd5
; 
32'd32166: dataIn1 = 32'd6
; 
32'd32167: dataIn1 = 32'd7
; 
32'd32168: dataIn1 = 32'd8
; 
32'd32169: dataIn1 = 32'd9
; 
32'd32170: dataIn1 = 32'd10
; 
32'd32171: dataIn1 = 32'd11
; 
32'd32172: dataIn1 = 32'd13
; 
32'd32173: dataIn1 = 32'd14
; 
32'd32174: dataIn1 = 32'd15
; 
32'd32175: dataIn1 = 32'd16
; 
32'd32176: dataIn1 = 32'd17
; 
32'd32177: dataIn1 = 32'd19
; 
32'd32178: dataIn1 = 32'd20
; 
32'd32179: dataIn1 = 32'd22
; 
32'd32180: dataIn1 = 32'd23
; 
32'd32181: dataIn1 = 32'd25
; 
32'd32182: dataIn1 = 32'd27
; 
32'd32183: dataIn1 = 32'd28
; 
32'd32184: dataIn1 = 32'd29
; 
32'd32185: dataIn1 = 32'd30
; 
32'd32186: dataIn1 = 32'd31
; 
32'd32187: dataIn1 = 32'd32
; 
32'd32188: dataIn1 = 32'd34
; 
32'd32189: dataIn1 = 32'd36
; 
32'd32190: dataIn1 = 32'd37
; 
32'd32191: dataIn1 = 32'd41
; 
32'd32192: dataIn1 = 32'd44
; 
32'd32193: dataIn1 = 32'd46
; 
32'd32194: dataIn1 = 32'd47
; 
32'd32195: dataIn1 = 32'd50
; 
32'd32196: dataIn1 = 32'd51
; 
32'd32197: dataIn1 = 32'd52
; 
32'd32198: dataIn1 = 32'd54
; 
32'd32199: dataIn1 = 32'd56
; 
32'd32200: dataIn1 = 32'd59
; 
32'd32201: dataIn1 = 32'd62
; 
32'd32202: dataIn1 = 32'd0
; 
32'd32203: dataIn1 = 32'd1
; 
32'd32204: dataIn1 = 32'd2
; 
32'd32205: dataIn1 = 32'd3
; 
32'd32206: dataIn1 = 32'd4
; 
32'd32207: dataIn1 = 32'd5
; 
32'd32208: dataIn1 = 32'd6
; 
32'd32209: dataIn1 = 32'd7
; 
32'd32210: dataIn1 = 32'd10
; 
32'd32211: dataIn1 = 32'd11
; 
32'd32212: dataIn1 = 32'd12
; 
32'd32213: dataIn1 = 32'd14
; 
32'd32214: dataIn1 = 32'd19
; 
32'd32215: dataIn1 = 32'd20
; 
32'd32216: dataIn1 = 32'd22
; 
32'd32217: dataIn1 = 32'd23
; 
32'd32218: dataIn1 = 32'd24
; 
32'd32219: dataIn1 = 32'd25
; 
32'd32220: dataIn1 = 32'd26
; 
32'd32221: dataIn1 = 32'd27
; 
32'd32222: dataIn1 = 32'd28
; 
32'd32223: dataIn1 = 32'd30
; 
32'd32224: dataIn1 = 32'd31
; 
32'd32225: dataIn1 = 32'd32
; 
32'd32226: dataIn1 = 32'd33
; 
32'd32227: dataIn1 = 32'd34
; 
32'd32228: dataIn1 = 32'd35
; 
32'd32229: dataIn1 = 32'd36
; 
32'd32230: dataIn1 = 32'd37
; 
32'd32231: dataIn1 = 32'd38
; 
32'd32232: dataIn1 = 32'd39
; 
32'd32233: dataIn1 = 32'd40
; 
32'd32234: dataIn1 = 32'd42
; 
32'd32235: dataIn1 = 32'd43
; 
32'd32236: dataIn1 = 32'd48
; 
32'd32237: dataIn1 = 32'd50
; 
32'd32238: dataIn1 = 32'd51
; 
32'd32239: dataIn1 = 32'd52
; 
32'd32240: dataIn1 = 32'd53
; 
32'd32241: dataIn1 = 32'd54
; 
32'd32242: dataIn1 = 32'd55
; 
32'd32243: dataIn1 = 32'd57
; 
32'd32244: dataIn1 = 32'd58
; 
32'd32245: dataIn1 = 32'd59
; 
32'd32246: dataIn1 = 32'd60
; 
32'd32247: dataIn1 = 32'd62
; 
32'd32248: dataIn1 = 32'd0
; 
32'd32249: dataIn1 = 32'd1
; 
32'd32250: dataIn1 = 32'd2
; 
32'd32251: dataIn1 = 32'd4
; 
32'd32252: dataIn1 = 32'd5
; 
32'd32253: dataIn1 = 32'd6
; 
32'd32254: dataIn1 = 32'd7
; 
32'd32255: dataIn1 = 32'd8
; 
32'd32256: dataIn1 = 32'd10
; 
32'd32257: dataIn1 = 32'd11
; 
32'd32258: dataIn1 = 32'd12
; 
32'd32259: dataIn1 = 32'd14
; 
32'd32260: dataIn1 = 32'd15
; 
32'd32261: dataIn1 = 32'd16
; 
32'd32262: dataIn1 = 32'd17
; 
32'd32263: dataIn1 = 32'd19
; 
32'd32264: dataIn1 = 32'd20
; 
32'd32265: dataIn1 = 32'd21
; 
32'd32266: dataIn1 = 32'd22
; 
32'd32267: dataIn1 = 32'd23
; 
32'd32268: dataIn1 = 32'd24
; 
32'd32269: dataIn1 = 32'd26
; 
32'd32270: dataIn1 = 32'd28
; 
32'd32271: dataIn1 = 32'd31
; 
32'd32272: dataIn1 = 32'd32
; 
32'd32273: dataIn1 = 32'd33
; 
32'd32274: dataIn1 = 32'd34
; 
32'd32275: dataIn1 = 32'd36
; 
32'd32276: dataIn1 = 32'd37
; 
32'd32277: dataIn1 = 32'd38
; 
32'd32278: dataIn1 = 32'd39
; 
32'd32279: dataIn1 = 32'd41
; 
32'd32280: dataIn1 = 32'd42
; 
32'd32281: dataIn1 = 32'd43
; 
32'd32282: dataIn1 = 32'd50
; 
32'd32283: dataIn1 = 32'd53
; 
32'd32284: dataIn1 = 32'd54
; 
32'd32285: dataIn1 = 32'd55
; 
32'd32286: dataIn1 = 32'd56
; 
32'd32287: dataIn1 = 32'd57
; 
32'd32288: dataIn1 = 32'd58
; 
32'd32289: dataIn1 = 32'd59
; 
32'd32290: dataIn1 = 32'd60
; 
32'd32291: dataIn1 = 32'd62
; 
32'd32292: dataIn1 = 32'd63
; 
32'd32293: dataIn1 = 32'd0
; 
32'd32294: dataIn1 = 32'd1
; 
32'd32295: dataIn1 = 32'd2
; 
32'd32296: dataIn1 = 32'd4
; 
32'd32297: dataIn1 = 32'd6
; 
32'd32298: dataIn1 = 32'd9
; 
32'd32299: dataIn1 = 32'd10
; 
32'd32300: dataIn1 = 32'd11
; 
32'd32301: dataIn1 = 32'd14
; 
32'd32302: dataIn1 = 32'd15
; 
32'd32303: dataIn1 = 32'd16
; 
32'd32304: dataIn1 = 32'd17
; 
32'd32305: dataIn1 = 32'd19
; 
32'd32306: dataIn1 = 32'd20
; 
32'd32307: dataIn1 = 32'd22
; 
32'd32308: dataIn1 = 32'd23
; 
32'd32309: dataIn1 = 32'd24
; 
32'd32310: dataIn1 = 32'd25
; 
32'd32311: dataIn1 = 32'd27
; 
32'd32312: dataIn1 = 32'd28
; 
32'd32313: dataIn1 = 32'd29
; 
32'd32314: dataIn1 = 32'd32
; 
32'd32315: dataIn1 = 32'd34
; 
32'd32316: dataIn1 = 32'd36
; 
32'd32317: dataIn1 = 32'd37
; 
32'd32318: dataIn1 = 32'd38
; 
32'd32319: dataIn1 = 32'd39
; 
32'd32320: dataIn1 = 32'd41
; 
32'd32321: dataIn1 = 32'd42
; 
32'd32322: dataIn1 = 32'd43
; 
32'd32323: dataIn1 = 32'd45
; 
32'd32324: dataIn1 = 32'd46
; 
32'd32325: dataIn1 = 32'd48
; 
32'd32326: dataIn1 = 32'd50
; 
32'd32327: dataIn1 = 32'd51
; 
32'd32328: dataIn1 = 32'd53
; 
32'd32329: dataIn1 = 32'd56
; 
32'd32330: dataIn1 = 32'd57
; 
32'd32331: dataIn1 = 32'd58
; 
32'd32332: dataIn1 = 32'd59
; 
32'd32333: dataIn1 = 32'd60
; 
32'd32334: dataIn1 = 32'd61
; 
32'd32335: dataIn1 = 32'd63
; 
32'd32336: dataIn1 = 32'd0
; 
32'd32337: dataIn1 = 32'd3
; 
32'd32338: dataIn1 = 32'd5
; 
32'd32339: dataIn1 = 32'd6
; 
32'd32340: dataIn1 = 32'd7
; 
32'd32341: dataIn1 = 32'd9
; 
32'd32342: dataIn1 = 32'd10
; 
32'd32343: dataIn1 = 32'd11
; 
32'd32344: dataIn1 = 32'd12
; 
32'd32345: dataIn1 = 32'd13
; 
32'd32346: dataIn1 = 32'd14
; 
32'd32347: dataIn1 = 32'd15
; 
32'd32348: dataIn1 = 32'd16
; 
32'd32349: dataIn1 = 32'd17
; 
32'd32350: dataIn1 = 32'd19
; 
32'd32351: dataIn1 = 32'd20
; 
32'd32352: dataIn1 = 32'd21
; 
32'd32353: dataIn1 = 32'd22
; 
32'd32354: dataIn1 = 32'd23
; 
32'd32355: dataIn1 = 32'd24
; 
32'd32356: dataIn1 = 32'd26
; 
32'd32357: dataIn1 = 32'd27
; 
32'd32358: dataIn1 = 32'd28
; 
32'd32359: dataIn1 = 32'd30
; 
32'd32360: dataIn1 = 32'd31
; 
32'd32361: dataIn1 = 32'd33
; 
32'd32362: dataIn1 = 32'd34
; 
32'd32363: dataIn1 = 32'd35
; 
32'd32364: dataIn1 = 32'd36
; 
32'd32365: dataIn1 = 32'd37
; 
32'd32366: dataIn1 = 32'd38
; 
32'd32367: dataIn1 = 32'd41
; 
32'd32368: dataIn1 = 32'd42
; 
32'd32369: dataIn1 = 32'd43
; 
32'd32370: dataIn1 = 32'd44
; 
32'd32371: dataIn1 = 32'd47
; 
32'd32372: dataIn1 = 32'd48
; 
32'd32373: dataIn1 = 32'd49
; 
32'd32374: dataIn1 = 32'd50
; 
32'd32375: dataIn1 = 32'd51
; 
32'd32376: dataIn1 = 32'd52
; 
32'd32377: dataIn1 = 32'd54
; 
32'd32378: dataIn1 = 32'd56
; 
32'd32379: dataIn1 = 32'd57
; 
32'd32380: dataIn1 = 32'd58
; 
32'd32381: dataIn1 = 32'd59
; 
32'd32382: dataIn1 = 32'd61
; 
32'd32383: dataIn1 = 32'd62
; 
32'd32384: dataIn1 = 32'd63
; 
32'd32385: dataIn1 = 32'd0
; 
32'd32386: dataIn1 = 32'd4
; 
32'd32387: dataIn1 = 32'd6
; 
32'd32388: dataIn1 = 32'd10
; 
32'd32389: dataIn1 = 32'd12
; 
32'd32390: dataIn1 = 32'd15
; 
32'd32391: dataIn1 = 32'd16
; 
32'd32392: dataIn1 = 32'd17
; 
32'd32393: dataIn1 = 32'd19
; 
32'd32394: dataIn1 = 32'd21
; 
32'd32395: dataIn1 = 32'd24
; 
32'd32396: dataIn1 = 32'd26
; 
32'd32397: dataIn1 = 32'd27
; 
32'd32398: dataIn1 = 32'd28
; 
32'd32399: dataIn1 = 32'd32
; 
32'd32400: dataIn1 = 32'd33
; 
32'd32401: dataIn1 = 32'd38
; 
32'd32402: dataIn1 = 32'd39
; 
32'd32403: dataIn1 = 32'd40
; 
32'd32404: dataIn1 = 32'd41
; 
32'd32405: dataIn1 = 32'd46
; 
32'd32406: dataIn1 = 32'd47
; 
32'd32407: dataIn1 = 32'd48
; 
32'd32408: dataIn1 = 32'd49
; 
32'd32409: dataIn1 = 32'd50
; 
32'd32410: dataIn1 = 32'd51
; 
32'd32411: dataIn1 = 32'd52
; 
32'd32412: dataIn1 = 32'd53
; 
32'd32413: dataIn1 = 32'd54
; 
32'd32414: dataIn1 = 32'd55
; 
32'd32415: dataIn1 = 32'd56
; 
32'd32416: dataIn1 = 32'd57
; 
32'd32417: dataIn1 = 32'd58
; 
32'd32418: dataIn1 = 32'd60
; 
32'd32419: dataIn1 = 32'd61
; 
32'd32420: dataIn1 = 32'd0
; 
32'd32421: dataIn1 = 32'd1
; 
32'd32422: dataIn1 = 32'd2
; 
32'd32423: dataIn1 = 32'd4
; 
32'd32424: dataIn1 = 32'd5
; 
32'd32425: dataIn1 = 32'd6
; 
32'd32426: dataIn1 = 32'd7
; 
32'd32427: dataIn1 = 32'd8
; 
32'd32428: dataIn1 = 32'd9
; 
32'd32429: dataIn1 = 32'd11
; 
32'd32430: dataIn1 = 32'd13
; 
32'd32431: dataIn1 = 32'd14
; 
32'd32432: dataIn1 = 32'd15
; 
32'd32433: dataIn1 = 32'd19
; 
32'd32434: dataIn1 = 32'd20
; 
32'd32435: dataIn1 = 32'd21
; 
32'd32436: dataIn1 = 32'd22
; 
32'd32437: dataIn1 = 32'd23
; 
32'd32438: dataIn1 = 32'd26
; 
32'd32439: dataIn1 = 32'd27
; 
32'd32440: dataIn1 = 32'd28
; 
32'd32441: dataIn1 = 32'd29
; 
32'd32442: dataIn1 = 32'd31
; 
32'd32443: dataIn1 = 32'd33
; 
32'd32444: dataIn1 = 32'd34
; 
32'd32445: dataIn1 = 32'd35
; 
32'd32446: dataIn1 = 32'd36
; 
32'd32447: dataIn1 = 32'd37
; 
32'd32448: dataIn1 = 32'd38
; 
32'd32449: dataIn1 = 32'd39
; 
32'd32450: dataIn1 = 32'd41
; 
32'd32451: dataIn1 = 32'd42
; 
32'd32452: dataIn1 = 32'd43
; 
32'd32453: dataIn1 = 32'd46
; 
32'd32454: dataIn1 = 32'd47
; 
32'd32455: dataIn1 = 32'd48
; 
32'd32456: dataIn1 = 32'd50
; 
32'd32457: dataIn1 = 32'd51
; 
32'd32458: dataIn1 = 32'd52
; 
32'd32459: dataIn1 = 32'd54
; 
32'd32460: dataIn1 = 32'd55
; 
32'd32461: dataIn1 = 32'd56
; 
32'd32462: dataIn1 = 32'd57
; 
32'd32463: dataIn1 = 32'd59
; 
32'd32464: dataIn1 = 32'd61
; 
32'd32465: dataIn1 = 32'd62
; 
32'd32466: dataIn1 = 32'd63
; 
32'd32467: dataIn1 = 32'd3
; 
32'd32468: dataIn1 = 32'd4
; 
32'd32469: dataIn1 = 32'd5
; 
32'd32470: dataIn1 = 32'd6
; 
32'd32471: dataIn1 = 32'd7
; 
32'd32472: dataIn1 = 32'd8
; 
32'd32473: dataIn1 = 32'd9
; 
32'd32474: dataIn1 = 32'd11
; 
32'd32475: dataIn1 = 32'd12
; 
32'd32476: dataIn1 = 32'd13
; 
32'd32477: dataIn1 = 32'd15
; 
32'd32478: dataIn1 = 32'd16
; 
32'd32479: dataIn1 = 32'd18
; 
32'd32480: dataIn1 = 32'd19
; 
32'd32481: dataIn1 = 32'd20
; 
32'd32482: dataIn1 = 32'd21
; 
32'd32483: dataIn1 = 32'd22
; 
32'd32484: dataIn1 = 32'd23
; 
32'd32485: dataIn1 = 32'd24
; 
32'd32486: dataIn1 = 32'd26
; 
32'd32487: dataIn1 = 32'd28
; 
32'd32488: dataIn1 = 32'd29
; 
32'd32489: dataIn1 = 32'd30
; 
32'd32490: dataIn1 = 32'd31
; 
32'd32491: dataIn1 = 32'd33
; 
32'd32492: dataIn1 = 32'd34
; 
32'd32493: dataIn1 = 32'd35
; 
32'd32494: dataIn1 = 32'd36
; 
32'd32495: dataIn1 = 32'd37
; 
32'd32496: dataIn1 = 32'd38
; 
32'd32497: dataIn1 = 32'd39
; 
32'd32498: dataIn1 = 32'd40
; 
32'd32499: dataIn1 = 32'd42
; 
32'd32500: dataIn1 = 32'd43
; 
32'd32501: dataIn1 = 32'd45
; 
32'd32502: dataIn1 = 32'd46
; 
32'd32503: dataIn1 = 32'd47
; 
32'd32504: dataIn1 = 32'd48
; 
32'd32505: dataIn1 = 32'd49
; 
32'd32506: dataIn1 = 32'd50
; 
32'd32507: dataIn1 = 32'd51
; 
32'd32508: dataIn1 = 32'd52
; 
32'd32509: dataIn1 = 32'd53
; 
32'd32510: dataIn1 = 32'd54
; 
32'd32511: dataIn1 = 32'd55
; 
32'd32512: dataIn1 = 32'd56
; 
32'd32513: dataIn1 = 32'd57
; 
32'd32514: dataIn1 = 32'd58
; 
32'd32515: dataIn1 = 32'd60
; 
32'd32516: dataIn1 = 32'd63
; 
32'd32517: dataIn1 = 32'd2
; 
32'd32518: dataIn1 = 32'd3
; 
32'd32519: dataIn1 = 32'd5
; 
32'd32520: dataIn1 = 32'd6
; 
32'd32521: dataIn1 = 32'd7
; 
32'd32522: dataIn1 = 32'd9
; 
32'd32523: dataIn1 = 32'd10
; 
32'd32524: dataIn1 = 32'd12
; 
32'd32525: dataIn1 = 32'd13
; 
32'd32526: dataIn1 = 32'd15
; 
32'd32527: dataIn1 = 32'd16
; 
32'd32528: dataIn1 = 32'd17
; 
32'd32529: dataIn1 = 32'd19
; 
32'd32530: dataIn1 = 32'd20
; 
32'd32531: dataIn1 = 32'd23
; 
32'd32532: dataIn1 = 32'd24
; 
32'd32533: dataIn1 = 32'd25
; 
32'd32534: dataIn1 = 32'd26
; 
32'd32535: dataIn1 = 32'd27
; 
32'd32536: dataIn1 = 32'd28
; 
32'd32537: dataIn1 = 32'd29
; 
32'd32538: dataIn1 = 32'd30
; 
32'd32539: dataIn1 = 32'd33
; 
32'd32540: dataIn1 = 32'd34
; 
32'd32541: dataIn1 = 32'd37
; 
32'd32542: dataIn1 = 32'd40
; 
32'd32543: dataIn1 = 32'd41
; 
32'd32544: dataIn1 = 32'd44
; 
32'd32545: dataIn1 = 32'd46
; 
32'd32546: dataIn1 = 32'd47
; 
32'd32547: dataIn1 = 32'd48
; 
32'd32548: dataIn1 = 32'd50
; 
32'd32549: dataIn1 = 32'd51
; 
32'd32550: dataIn1 = 32'd52
; 
32'd32551: dataIn1 = 32'd55
; 
32'd32552: dataIn1 = 32'd56
; 
32'd32553: dataIn1 = 32'd57
; 
32'd32554: dataIn1 = 32'd58
; 
32'd32555: dataIn1 = 32'd60
; 
32'd32556: dataIn1 = 32'd61
; 
32'd32557: dataIn1 = 32'd62
; 
32'd32558: dataIn1 = 32'd63
; 
32'd32559: dataIn1 = 32'd1
; 
32'd32560: dataIn1 = 32'd2
; 
32'd32561: dataIn1 = 32'd3
; 
32'd32562: dataIn1 = 32'd7
; 
32'd32563: dataIn1 = 32'd8
; 
32'd32564: dataIn1 = 32'd9
; 
32'd32565: dataIn1 = 32'd10
; 
32'd32566: dataIn1 = 32'd11
; 
32'd32567: dataIn1 = 32'd13
; 
32'd32568: dataIn1 = 32'd14
; 
32'd32569: dataIn1 = 32'd17
; 
32'd32570: dataIn1 = 32'd18
; 
32'd32571: dataIn1 = 32'd19
; 
32'd32572: dataIn1 = 32'd20
; 
32'd32573: dataIn1 = 32'd21
; 
32'd32574: dataIn1 = 32'd22
; 
32'd32575: dataIn1 = 32'd23
; 
32'd32576: dataIn1 = 32'd26
; 
32'd32577: dataIn1 = 32'd28
; 
32'd32578: dataIn1 = 32'd29
; 
32'd32579: dataIn1 = 32'd30
; 
32'd32580: dataIn1 = 32'd32
; 
32'd32581: dataIn1 = 32'd33
; 
32'd32582: dataIn1 = 32'd35
; 
32'd32583: dataIn1 = 32'd36
; 
32'd32584: dataIn1 = 32'd38
; 
32'd32585: dataIn1 = 32'd39
; 
32'd32586: dataIn1 = 32'd42
; 
32'd32587: dataIn1 = 32'd47
; 
32'd32588: dataIn1 = 32'd48
; 
32'd32589: dataIn1 = 32'd49
; 
32'd32590: dataIn1 = 32'd50
; 
32'd32591: dataIn1 = 32'd52
; 
32'd32592: dataIn1 = 32'd53
; 
32'd32593: dataIn1 = 32'd55
; 
32'd32594: dataIn1 = 32'd56
; 
32'd32595: dataIn1 = 32'd57
; 
32'd32596: dataIn1 = 32'd58
; 
32'd32597: dataIn1 = 32'd59
; 
32'd32598: dataIn1 = 32'd62
; 
32'd32599: dataIn1 = 32'd63
; 
32'd32600: dataIn1 = 32'd0
; 
32'd32601: dataIn1 = 32'd1
; 
32'd32602: dataIn1 = 32'd2
; 
32'd32603: dataIn1 = 32'd4
; 
32'd32604: dataIn1 = 32'd5
; 
32'd32605: dataIn1 = 32'd6
; 
32'd32606: dataIn1 = 32'd9
; 
32'd32607: dataIn1 = 32'd10
; 
32'd32608: dataIn1 = 32'd13
; 
32'd32609: dataIn1 = 32'd15
; 
32'd32610: dataIn1 = 32'd18
; 
32'd32611: dataIn1 = 32'd19
; 
32'd32612: dataIn1 = 32'd20
; 
32'd32613: dataIn1 = 32'd22
; 
32'd32614: dataIn1 = 32'd23
; 
32'd32615: dataIn1 = 32'd24
; 
32'd32616: dataIn1 = 32'd26
; 
32'd32617: dataIn1 = 32'd27
; 
32'd32618: dataIn1 = 32'd28
; 
32'd32619: dataIn1 = 32'd30
; 
32'd32620: dataIn1 = 32'd31
; 
32'd32621: dataIn1 = 32'd32
; 
32'd32622: dataIn1 = 32'd34
; 
32'd32623: dataIn1 = 32'd37
; 
32'd32624: dataIn1 = 32'd40
; 
32'd32625: dataIn1 = 32'd41
; 
32'd32626: dataIn1 = 32'd43
; 
32'd32627: dataIn1 = 32'd44
; 
32'd32628: dataIn1 = 32'd45
; 
32'd32629: dataIn1 = 32'd50
; 
32'd32630: dataIn1 = 32'd51
; 
32'd32631: dataIn1 = 32'd52
; 
32'd32632: dataIn1 = 32'd53
; 
32'd32633: dataIn1 = 32'd54
; 
32'd32634: dataIn1 = 32'd55
; 
32'd32635: dataIn1 = 32'd57
; 
32'd32636: dataIn1 = 32'd58
; 
32'd32637: dataIn1 = 32'd60
; 
32'd32638: dataIn1 = 32'd61
; 
32'd32639: dataIn1 = 32'd62
; 
32'd32640: dataIn1 = 32'd0
; 
32'd32641: dataIn1 = 32'd1
; 
32'd32642: dataIn1 = 32'd2
; 
32'd32643: dataIn1 = 32'd3
; 
32'd32644: dataIn1 = 32'd6
; 
32'd32645: dataIn1 = 32'd7
; 
32'd32646: dataIn1 = 32'd9
; 
32'd32647: dataIn1 = 32'd11
; 
32'd32648: dataIn1 = 32'd12
; 
32'd32649: dataIn1 = 32'd13
; 
32'd32650: dataIn1 = 32'd14
; 
32'd32651: dataIn1 = 32'd15
; 
32'd32652: dataIn1 = 32'd18
; 
32'd32653: dataIn1 = 32'd19
; 
32'd32654: dataIn1 = 32'd20
; 
32'd32655: dataIn1 = 32'd23
; 
32'd32656: dataIn1 = 32'd25
; 
32'd32657: dataIn1 = 32'd26
; 
32'd32658: dataIn1 = 32'd28
; 
32'd32659: dataIn1 = 32'd30
; 
32'd32660: dataIn1 = 32'd32
; 
32'd32661: dataIn1 = 32'd35
; 
32'd32662: dataIn1 = 32'd37
; 
32'd32663: dataIn1 = 32'd38
; 
32'd32664: dataIn1 = 32'd39
; 
32'd32665: dataIn1 = 32'd40
; 
32'd32666: dataIn1 = 32'd41
; 
32'd32667: dataIn1 = 32'd42
; 
32'd32668: dataIn1 = 32'd43
; 
32'd32669: dataIn1 = 32'd44
; 
32'd32670: dataIn1 = 32'd45
; 
32'd32671: dataIn1 = 32'd46
; 
32'd32672: dataIn1 = 32'd47
; 
32'd32673: dataIn1 = 32'd49
; 
32'd32674: dataIn1 = 32'd51
; 
32'd32675: dataIn1 = 32'd52
; 
32'd32676: dataIn1 = 32'd53
; 
32'd32677: dataIn1 = 32'd54
; 
32'd32678: dataIn1 = 32'd55
; 
32'd32679: dataIn1 = 32'd56
; 
32'd32680: dataIn1 = 32'd57
; 
32'd32681: dataIn1 = 32'd58
; 
32'd32682: dataIn1 = 32'd59
; 
32'd32683: dataIn1 = 32'd60
; 
32'd32684: dataIn1 = 32'd62
; 
32'd32685: dataIn1 = 32'd1
; 
32'd32686: dataIn1 = 32'd2
; 
32'd32687: dataIn1 = 32'd4
; 
32'd32688: dataIn1 = 32'd5
; 
32'd32689: dataIn1 = 32'd8
; 
32'd32690: dataIn1 = 32'd11
; 
32'd32691: dataIn1 = 32'd15
; 
32'd32692: dataIn1 = 32'd17
; 
32'd32693: dataIn1 = 32'd18
; 
32'd32694: dataIn1 = 32'd19
; 
32'd32695: dataIn1 = 32'd20
; 
32'd32696: dataIn1 = 32'd21
; 
32'd32697: dataIn1 = 32'd22
; 
32'd32698: dataIn1 = 32'd23
; 
32'd32699: dataIn1 = 32'd25
; 
32'd32700: dataIn1 = 32'd26
; 
32'd32701: dataIn1 = 32'd27
; 
32'd32702: dataIn1 = 32'd28
; 
32'd32703: dataIn1 = 32'd29
; 
32'd32704: dataIn1 = 32'd30
; 
32'd32705: dataIn1 = 32'd31
; 
32'd32706: dataIn1 = 32'd32
; 
32'd32707: dataIn1 = 32'd34
; 
32'd32708: dataIn1 = 32'd35
; 
32'd32709: dataIn1 = 32'd39
; 
32'd32710: dataIn1 = 32'd40
; 
32'd32711: dataIn1 = 32'd42
; 
32'd32712: dataIn1 = 32'd44
; 
32'd32713: dataIn1 = 32'd45
; 
32'd32714: dataIn1 = 32'd46
; 
32'd32715: dataIn1 = 32'd47
; 
32'd32716: dataIn1 = 32'd48
; 
32'd32717: dataIn1 = 32'd50
; 
32'd32718: dataIn1 = 32'd51
; 
32'd32719: dataIn1 = 32'd52
; 
32'd32720: dataIn1 = 32'd53
; 
32'd32721: dataIn1 = 32'd54
; 
32'd32722: dataIn1 = 32'd55
; 
32'd32723: dataIn1 = 32'd57
; 
32'd32724: dataIn1 = 32'd62
; 
32'd32725: dataIn1 = 32'd63
; 
32'd32726: dataIn1 = 32'd0
; 
32'd32727: dataIn1 = 32'd1
; 
32'd32728: dataIn1 = 32'd2
; 
32'd32729: dataIn1 = 32'd3
; 
32'd32730: dataIn1 = 32'd4
; 
32'd32731: dataIn1 = 32'd5
; 
32'd32732: dataIn1 = 32'd6
; 
32'd32733: dataIn1 = 32'd7
; 
32'd32734: dataIn1 = 32'd8
; 
32'd32735: dataIn1 = 32'd10
; 
32'd32736: dataIn1 = 32'd11
; 
32'd32737: dataIn1 = 32'd12
; 
32'd32738: dataIn1 = 32'd13
; 
32'd32739: dataIn1 = 32'd14
; 
32'd32740: dataIn1 = 32'd15
; 
32'd32741: dataIn1 = 32'd16
; 
32'd32742: dataIn1 = 32'd17
; 
32'd32743: dataIn1 = 32'd19
; 
32'd32744: dataIn1 = 32'd20
; 
32'd32745: dataIn1 = 32'd21
; 
32'd32746: dataIn1 = 32'd22
; 
32'd32747: dataIn1 = 32'd23
; 
32'd32748: dataIn1 = 32'd24
; 
32'd32749: dataIn1 = 32'd26
; 
32'd32750: dataIn1 = 32'd29
; 
32'd32751: dataIn1 = 32'd33
; 
32'd32752: dataIn1 = 32'd34
; 
32'd32753: dataIn1 = 32'd35
; 
32'd32754: dataIn1 = 32'd39
; 
32'd32755: dataIn1 = 32'd40
; 
32'd32756: dataIn1 = 32'd41
; 
32'd32757: dataIn1 = 32'd42
; 
32'd32758: dataIn1 = 32'd43
; 
32'd32759: dataIn1 = 32'd44
; 
32'd32760: dataIn1 = 32'd45
; 
32'd32761: dataIn1 = 32'd46
; 
32'd32762: dataIn1 = 32'd47
; 
32'd32763: dataIn1 = 32'd48
; 
32'd32764: dataIn1 = 32'd49
; 
32'd32765: dataIn1 = 32'd50
; 
32'd32766: dataIn1 = 32'd51
; 
32'd32767: dataIn1 = 32'd52
; 
32'd32768: dataIn1 = 32'd53
; 
32'd32769: dataIn1 = 32'd54
; 
32'd32770: dataIn1 = 32'd55
; 
32'd32771: dataIn1 = 32'd56
; 
32'd32772: dataIn1 = 32'd57
; 
32'd32773: dataIn1 = 32'd60
; 
32'd32774: dataIn1 = 32'd61
; 
32'd32775: dataIn1 = 32'd62
; 
32'd32776: dataIn1 = 32'd63
; 
32'd32777: dataIn1 = 32'd1
; 
32'd32778: dataIn1 = 32'd2
; 
32'd32779: dataIn1 = 32'd3
; 
32'd32780: dataIn1 = 32'd4
; 
32'd32781: dataIn1 = 32'd5
; 
32'd32782: dataIn1 = 32'd6
; 
32'd32783: dataIn1 = 32'd7
; 
32'd32784: dataIn1 = 32'd11
; 
32'd32785: dataIn1 = 32'd13
; 
32'd32786: dataIn1 = 32'd14
; 
32'd32787: dataIn1 = 32'd15
; 
32'd32788: dataIn1 = 32'd16
; 
32'd32789: dataIn1 = 32'd19
; 
32'd32790: dataIn1 = 32'd20
; 
32'd32791: dataIn1 = 32'd24
; 
32'd32792: dataIn1 = 32'd26
; 
32'd32793: dataIn1 = 32'd27
; 
32'd32794: dataIn1 = 32'd29
; 
32'd32795: dataIn1 = 32'd30
; 
32'd32796: dataIn1 = 32'd32
; 
32'd32797: dataIn1 = 32'd33
; 
32'd32798: dataIn1 = 32'd34
; 
32'd32799: dataIn1 = 32'd35
; 
32'd32800: dataIn1 = 32'd36
; 
32'd32801: dataIn1 = 32'd37
; 
32'd32802: dataIn1 = 32'd39
; 
32'd32803: dataIn1 = 32'd40
; 
32'd32804: dataIn1 = 32'd41
; 
32'd32805: dataIn1 = 32'd43
; 
32'd32806: dataIn1 = 32'd45
; 
32'd32807: dataIn1 = 32'd47
; 
32'd32808: dataIn1 = 32'd48
; 
32'd32809: dataIn1 = 32'd49
; 
32'd32810: dataIn1 = 32'd52
; 
32'd32811: dataIn1 = 32'd56
; 
32'd32812: dataIn1 = 32'd57
; 
32'd32813: dataIn1 = 32'd58
; 
32'd32814: dataIn1 = 32'd60
; 
32'd32815: dataIn1 = 32'd62
; 
32'd32816: dataIn1 = 32'd63
; 
32'd32817: dataIn1 = 32'd0
; 
32'd32818: dataIn1 = 32'd1
; 
32'd32819: dataIn1 = 32'd2
; 
32'd32820: dataIn1 = 32'd3
; 
32'd32821: dataIn1 = 32'd7
; 
32'd32822: dataIn1 = 32'd8
; 
32'd32823: dataIn1 = 32'd9
; 
32'd32824: dataIn1 = 32'd10
; 
32'd32825: dataIn1 = 32'd11
; 
32'd32826: dataIn1 = 32'd12
; 
32'd32827: dataIn1 = 32'd13
; 
32'd32828: dataIn1 = 32'd17
; 
32'd32829: dataIn1 = 32'd18
; 
32'd32830: dataIn1 = 32'd21
; 
32'd32831: dataIn1 = 32'd23
; 
32'd32832: dataIn1 = 32'd24
; 
32'd32833: dataIn1 = 32'd25
; 
32'd32834: dataIn1 = 32'd26
; 
32'd32835: dataIn1 = 32'd27
; 
32'd32836: dataIn1 = 32'd28
; 
32'd32837: dataIn1 = 32'd29
; 
32'd32838: dataIn1 = 32'd31
; 
32'd32839: dataIn1 = 32'd32
; 
32'd32840: dataIn1 = 32'd33
; 
32'd32841: dataIn1 = 32'd35
; 
32'd32842: dataIn1 = 32'd36
; 
32'd32843: dataIn1 = 32'd37
; 
32'd32844: dataIn1 = 32'd38
; 
32'd32845: dataIn1 = 32'd40
; 
32'd32846: dataIn1 = 32'd42
; 
32'd32847: dataIn1 = 32'd43
; 
32'd32848: dataIn1 = 32'd44
; 
32'd32849: dataIn1 = 32'd45
; 
32'd32850: dataIn1 = 32'd47
; 
32'd32851: dataIn1 = 32'd48
; 
32'd32852: dataIn1 = 32'd49
; 
32'd32853: dataIn1 = 32'd50
; 
32'd32854: dataIn1 = 32'd51
; 
32'd32855: dataIn1 = 32'd52
; 
32'd32856: dataIn1 = 32'd54
; 
32'd32857: dataIn1 = 32'd55
; 
32'd32858: dataIn1 = 32'd56
; 
32'd32859: dataIn1 = 32'd57
; 
32'd32860: dataIn1 = 32'd60
; 
32'd32861: dataIn1 = 32'd0
; 
32'd32862: dataIn1 = 32'd1
; 
32'd32863: dataIn1 = 32'd2
; 
32'd32864: dataIn1 = 32'd4
; 
32'd32865: dataIn1 = 32'd5
; 
32'd32866: dataIn1 = 32'd6
; 
32'd32867: dataIn1 = 32'd7
; 
32'd32868: dataIn1 = 32'd9
; 
32'd32869: dataIn1 = 32'd10
; 
32'd32870: dataIn1 = 32'd11
; 
32'd32871: dataIn1 = 32'd12
; 
32'd32872: dataIn1 = 32'd13
; 
32'd32873: dataIn1 = 32'd14
; 
32'd32874: dataIn1 = 32'd15
; 
32'd32875: dataIn1 = 32'd16
; 
32'd32876: dataIn1 = 32'd17
; 
32'd32877: dataIn1 = 32'd18
; 
32'd32878: dataIn1 = 32'd19
; 
32'd32879: dataIn1 = 32'd20
; 
32'd32880: dataIn1 = 32'd21
; 
32'd32881: dataIn1 = 32'd22
; 
32'd32882: dataIn1 = 32'd25
; 
32'd32883: dataIn1 = 32'd26
; 
32'd32884: dataIn1 = 32'd28
; 
32'd32885: dataIn1 = 32'd31
; 
32'd32886: dataIn1 = 32'd32
; 
32'd32887: dataIn1 = 32'd34
; 
32'd32888: dataIn1 = 32'd35
; 
32'd32889: dataIn1 = 32'd36
; 
32'd32890: dataIn1 = 32'd38
; 
32'd32891: dataIn1 = 32'd39
; 
32'd32892: dataIn1 = 32'd40
; 
32'd32893: dataIn1 = 32'd41
; 
32'd32894: dataIn1 = 32'd42
; 
32'd32895: dataIn1 = 32'd43
; 
32'd32896: dataIn1 = 32'd44
; 
32'd32897: dataIn1 = 32'd47
; 
32'd32898: dataIn1 = 32'd50
; 
32'd32899: dataIn1 = 32'd51
; 
32'd32900: dataIn1 = 32'd52
; 
32'd32901: dataIn1 = 32'd53
; 
32'd32902: dataIn1 = 32'd56
; 
32'd32903: dataIn1 = 32'd58
; 
32'd32904: dataIn1 = 32'd59
; 
32'd32905: dataIn1 = 32'd60
; 
32'd32906: dataIn1 = 32'd61
; 
32'd32907: dataIn1 = 32'd62
; 
32'd32908: dataIn1 = 32'd63
; 
32'd32909: dataIn1 = 32'd0
; 
32'd32910: dataIn1 = 32'd1
; 
32'd32911: dataIn1 = 32'd4
; 
32'd32912: dataIn1 = 32'd5
; 
32'd32913: dataIn1 = 32'd6
; 
32'd32914: dataIn1 = 32'd8
; 
32'd32915: dataIn1 = 32'd9
; 
32'd32916: dataIn1 = 32'd12
; 
32'd32917: dataIn1 = 32'd15
; 
32'd32918: dataIn1 = 32'd16
; 
32'd32919: dataIn1 = 32'd17
; 
32'd32920: dataIn1 = 32'd20
; 
32'd32921: dataIn1 = 32'd21
; 
32'd32922: dataIn1 = 32'd24
; 
32'd32923: dataIn1 = 32'd25
; 
32'd32924: dataIn1 = 32'd26
; 
32'd32925: dataIn1 = 32'd27
; 
32'd32926: dataIn1 = 32'd29
; 
32'd32927: dataIn1 = 32'd31
; 
32'd32928: dataIn1 = 32'd34
; 
32'd32929: dataIn1 = 32'd35
; 
32'd32930: dataIn1 = 32'd37
; 
32'd32931: dataIn1 = 32'd39
; 
32'd32932: dataIn1 = 32'd40
; 
32'd32933: dataIn1 = 32'd41
; 
32'd32934: dataIn1 = 32'd42
; 
32'd32935: dataIn1 = 32'd43
; 
32'd32936: dataIn1 = 32'd46
; 
32'd32937: dataIn1 = 32'd47
; 
32'd32938: dataIn1 = 32'd48
; 
32'd32939: dataIn1 = 32'd49
; 
32'd32940: dataIn1 = 32'd50
; 
32'd32941: dataIn1 = 32'd52
; 
32'd32942: dataIn1 = 32'd55
; 
32'd32943: dataIn1 = 32'd56
; 
32'd32944: dataIn1 = 32'd57
; 
32'd32945: dataIn1 = 32'd58
; 
32'd32946: dataIn1 = 32'd59
; 
32'd32947: dataIn1 = 32'd60
; 
32'd32948: dataIn1 = 32'd61
; 
32'd32949: dataIn1 = 32'd62
; 
32'd32950: dataIn1 = 32'd63
; 
32'd32951: dataIn1 = 32'd0
; 
32'd32952: dataIn1 = 32'd1
; 
32'd32953: dataIn1 = 32'd2
; 
32'd32954: dataIn1 = 32'd3
; 
32'd32955: dataIn1 = 32'd4
; 
32'd32956: dataIn1 = 32'd7
; 
32'd32957: dataIn1 = 32'd8
; 
32'd32958: dataIn1 = 32'd9
; 
32'd32959: dataIn1 = 32'd11
; 
32'd32960: dataIn1 = 32'd13
; 
32'd32961: dataIn1 = 32'd14
; 
32'd32962: dataIn1 = 32'd16
; 
32'd32963: dataIn1 = 32'd17
; 
32'd32964: dataIn1 = 32'd19
; 
32'd32965: dataIn1 = 32'd20
; 
32'd32966: dataIn1 = 32'd22
; 
32'd32967: dataIn1 = 32'd23
; 
32'd32968: dataIn1 = 32'd24
; 
32'd32969: dataIn1 = 32'd25
; 
32'd32970: dataIn1 = 32'd26
; 
32'd32971: dataIn1 = 32'd27
; 
32'd32972: dataIn1 = 32'd28
; 
32'd32973: dataIn1 = 32'd29
; 
32'd32974: dataIn1 = 32'd30
; 
32'd32975: dataIn1 = 32'd32
; 
32'd32976: dataIn1 = 32'd33
; 
32'd32977: dataIn1 = 32'd35
; 
32'd32978: dataIn1 = 32'd37
; 
32'd32979: dataIn1 = 32'd39
; 
32'd32980: dataIn1 = 32'd40
; 
32'd32981: dataIn1 = 32'd41
; 
32'd32982: dataIn1 = 32'd45
; 
32'd32983: dataIn1 = 32'd46
; 
32'd32984: dataIn1 = 32'd47
; 
32'd32985: dataIn1 = 32'd48
; 
32'd32986: dataIn1 = 32'd49
; 
32'd32987: dataIn1 = 32'd50
; 
32'd32988: dataIn1 = 32'd51
; 
32'd32989: dataIn1 = 32'd53
; 
32'd32990: dataIn1 = 32'd54
; 
32'd32991: dataIn1 = 32'd55
; 
32'd32992: dataIn1 = 32'd56
; 
32'd32993: dataIn1 = 32'd58
; 
32'd32994: dataIn1 = 32'd59
; 
32'd32995: dataIn1 = 32'd60
; 
32'd32996: dataIn1 = 32'd61
; 
32'd32997: dataIn1 = 32'd62
; 
32'd32998: dataIn1 = 32'd63
; 
32'd32999: dataIn1 = 32'd0
; 
32'd33000: dataIn1 = 32'd2
; 
32'd33001: dataIn1 = 32'd3
; 
32'd33002: dataIn1 = 32'd5
; 
32'd33003: dataIn1 = 32'd6
; 
32'd33004: dataIn1 = 32'd7
; 
32'd33005: dataIn1 = 32'd8
; 
32'd33006: dataIn1 = 32'd9
; 
32'd33007: dataIn1 = 32'd12
; 
32'd33008: dataIn1 = 32'd13
; 
32'd33009: dataIn1 = 32'd15
; 
32'd33010: dataIn1 = 32'd16
; 
32'd33011: dataIn1 = 32'd18
; 
32'd33012: dataIn1 = 32'd19
; 
32'd33013: dataIn1 = 32'd20
; 
32'd33014: dataIn1 = 32'd21
; 
32'd33015: dataIn1 = 32'd22
; 
32'd33016: dataIn1 = 32'd25
; 
32'd33017: dataIn1 = 32'd27
; 
32'd33018: dataIn1 = 32'd29
; 
32'd33019: dataIn1 = 32'd31
; 
32'd33020: dataIn1 = 32'd32
; 
32'd33021: dataIn1 = 32'd34
; 
32'd33022: dataIn1 = 32'd36
; 
32'd33023: dataIn1 = 32'd37
; 
32'd33024: dataIn1 = 32'd38
; 
32'd33025: dataIn1 = 32'd39
; 
32'd33026: dataIn1 = 32'd40
; 
32'd33027: dataIn1 = 32'd41
; 
32'd33028: dataIn1 = 32'd42
; 
32'd33029: dataIn1 = 32'd43
; 
32'd33030: dataIn1 = 32'd44
; 
32'd33031: dataIn1 = 32'd48
; 
32'd33032: dataIn1 = 32'd49
; 
32'd33033: dataIn1 = 32'd50
; 
32'd33034: dataIn1 = 32'd51
; 
32'd33035: dataIn1 = 32'd52
; 
32'd33036: dataIn1 = 32'd53
; 
32'd33037: dataIn1 = 32'd57
; 
32'd33038: dataIn1 = 32'd59
; 
32'd33039: dataIn1 = 32'd61
; 
32'd33040: dataIn1 = 32'd62
; 
32'd33041: dataIn1 = 32'd63
; 
32'd33042: dataIn1 = 32'd1
; 
32'd33043: dataIn1 = 32'd3
; 
32'd33044: dataIn1 = 32'd4
; 
32'd33045: dataIn1 = 32'd5
; 
32'd33046: dataIn1 = 32'd6
; 
32'd33047: dataIn1 = 32'd7
; 
32'd33048: dataIn1 = 32'd9
; 
32'd33049: dataIn1 = 32'd10
; 
32'd33050: dataIn1 = 32'd12
; 
32'd33051: dataIn1 = 32'd13
; 
32'd33052: dataIn1 = 32'd14
; 
32'd33053: dataIn1 = 32'd15
; 
32'd33054: dataIn1 = 32'd16
; 
32'd33055: dataIn1 = 32'd19
; 
32'd33056: dataIn1 = 32'd20
; 
32'd33057: dataIn1 = 32'd21
; 
32'd33058: dataIn1 = 32'd22
; 
32'd33059: dataIn1 = 32'd23
; 
32'd33060: dataIn1 = 32'd24
; 
32'd33061: dataIn1 = 32'd25
; 
32'd33062: dataIn1 = 32'd26
; 
32'd33063: dataIn1 = 32'd27
; 
32'd33064: dataIn1 = 32'd28
; 
32'd33065: dataIn1 = 32'd29
; 
32'd33066: dataIn1 = 32'd30
; 
32'd33067: dataIn1 = 32'd31
; 
32'd33068: dataIn1 = 32'd34
; 
32'd33069: dataIn1 = 32'd36
; 
32'd33070: dataIn1 = 32'd37
; 
32'd33071: dataIn1 = 32'd38
; 
32'd33072: dataIn1 = 32'd39
; 
32'd33073: dataIn1 = 32'd41
; 
32'd33074: dataIn1 = 32'd42
; 
32'd33075: dataIn1 = 32'd43
; 
32'd33076: dataIn1 = 32'd45
; 
32'd33077: dataIn1 = 32'd49
; 
32'd33078: dataIn1 = 32'd50
; 
32'd33079: dataIn1 = 32'd51
; 
32'd33080: dataIn1 = 32'd52
; 
32'd33081: dataIn1 = 32'd53
; 
32'd33082: dataIn1 = 32'd54
; 
32'd33083: dataIn1 = 32'd55
; 
32'd33084: dataIn1 = 32'd56
; 
32'd33085: dataIn1 = 32'd59
; 
32'd33086: dataIn1 = 32'd60
; 
32'd33087: dataIn1 = 32'd62
; 
32'd33088: dataIn1 = 32'd63
; 
32'd33089: dataIn1 = 32'd0
; 
32'd33090: dataIn1 = 32'd1
; 
32'd33091: dataIn1 = 32'd2
; 
32'd33092: dataIn1 = 32'd3
; 
32'd33093: dataIn1 = 32'd4
; 
32'd33094: dataIn1 = 32'd5
; 
32'd33095: dataIn1 = 32'd6
; 
32'd33096: dataIn1 = 32'd7
; 
32'd33097: dataIn1 = 32'd9
; 
32'd33098: dataIn1 = 32'd10
; 
32'd33099: dataIn1 = 32'd11
; 
32'd33100: dataIn1 = 32'd14
; 
32'd33101: dataIn1 = 32'd15
; 
32'd33102: dataIn1 = 32'd16
; 
32'd33103: dataIn1 = 32'd18
; 
32'd33104: dataIn1 = 32'd19
; 
32'd33105: dataIn1 = 32'd21
; 
32'd33106: dataIn1 = 32'd22
; 
32'd33107: dataIn1 = 32'd23
; 
32'd33108: dataIn1 = 32'd26
; 
32'd33109: dataIn1 = 32'd27
; 
32'd33110: dataIn1 = 32'd28
; 
32'd33111: dataIn1 = 32'd29
; 
32'd33112: dataIn1 = 32'd30
; 
32'd33113: dataIn1 = 32'd31
; 
32'd33114: dataIn1 = 32'd32
; 
32'd33115: dataIn1 = 32'd33
; 
32'd33116: dataIn1 = 32'd34
; 
32'd33117: dataIn1 = 32'd36
; 
32'd33118: dataIn1 = 32'd37
; 
32'd33119: dataIn1 = 32'd38
; 
32'd33120: dataIn1 = 32'd40
; 
32'd33121: dataIn1 = 32'd41
; 
32'd33122: dataIn1 = 32'd42
; 
32'd33123: dataIn1 = 32'd44
; 
32'd33124: dataIn1 = 32'd45
; 
32'd33125: dataIn1 = 32'd46
; 
32'd33126: dataIn1 = 32'd50
; 
32'd33127: dataIn1 = 32'd52
; 
32'd33128: dataIn1 = 32'd53
; 
32'd33129: dataIn1 = 32'd54
; 
32'd33130: dataIn1 = 32'd55
; 
32'd33131: dataIn1 = 32'd56
; 
32'd33132: dataIn1 = 32'd57
; 
32'd33133: dataIn1 = 32'd58
; 
32'd33134: dataIn1 = 32'd59
; 
32'd33135: dataIn1 = 32'd60
; 
32'd33136: dataIn1 = 32'd63
; 
32'd33137: dataIn1 = 32'd0
; 
32'd33138: dataIn1 = 32'd2
; 
32'd33139: dataIn1 = 32'd3
; 
32'd33140: dataIn1 = 32'd4
; 
32'd33141: dataIn1 = 32'd5
; 
32'd33142: dataIn1 = 32'd8
; 
32'd33143: dataIn1 = 32'd9
; 
32'd33144: dataIn1 = 32'd10
; 
32'd33145: dataIn1 = 32'd11
; 
32'd33146: dataIn1 = 32'd12
; 
32'd33147: dataIn1 = 32'd13
; 
32'd33148: dataIn1 = 32'd16
; 
32'd33149: dataIn1 = 32'd17
; 
32'd33150: dataIn1 = 32'd18
; 
32'd33151: dataIn1 = 32'd19
; 
32'd33152: dataIn1 = 32'd20
; 
32'd33153: dataIn1 = 32'd22
; 
32'd33154: dataIn1 = 32'd23
; 
32'd33155: dataIn1 = 32'd24
; 
32'd33156: dataIn1 = 32'd25
; 
32'd33157: dataIn1 = 32'd26
; 
32'd33158: dataIn1 = 32'd27
; 
32'd33159: dataIn1 = 32'd30
; 
32'd33160: dataIn1 = 32'd32
; 
32'd33161: dataIn1 = 32'd33
; 
32'd33162: dataIn1 = 32'd34
; 
32'd33163: dataIn1 = 32'd36
; 
32'd33164: dataIn1 = 32'd37
; 
32'd33165: dataIn1 = 32'd39
; 
32'd33166: dataIn1 = 32'd40
; 
32'd33167: dataIn1 = 32'd42
; 
32'd33168: dataIn1 = 32'd45
; 
32'd33169: dataIn1 = 32'd46
; 
32'd33170: dataIn1 = 32'd50
; 
32'd33171: dataIn1 = 32'd51
; 
32'd33172: dataIn1 = 32'd53
; 
32'd33173: dataIn1 = 32'd54
; 
32'd33174: dataIn1 = 32'd55
; 
32'd33175: dataIn1 = 32'd57
; 
32'd33176: dataIn1 = 32'd58
; 
32'd33177: dataIn1 = 32'd59
; 
32'd33178: dataIn1 = 32'd60
; 
32'd33179: dataIn1 = 32'd61
; 
32'd33180: dataIn1 = 32'd1
; 
32'd33181: dataIn1 = 32'd3
; 
32'd33182: dataIn1 = 32'd4
; 
32'd33183: dataIn1 = 32'd5
; 
32'd33184: dataIn1 = 32'd6
; 
32'd33185: dataIn1 = 32'd7
; 
32'd33186: dataIn1 = 32'd8
; 
32'd33187: dataIn1 = 32'd9
; 
32'd33188: dataIn1 = 32'd10
; 
32'd33189: dataIn1 = 32'd11
; 
32'd33190: dataIn1 = 32'd12
; 
32'd33191: dataIn1 = 32'd13
; 
32'd33192: dataIn1 = 32'd14
; 
32'd33193: dataIn1 = 32'd15
; 
32'd33194: dataIn1 = 32'd16
; 
32'd33195: dataIn1 = 32'd18
; 
32'd33196: dataIn1 = 32'd20
; 
32'd33197: dataIn1 = 32'd24
; 
32'd33198: dataIn1 = 32'd25
; 
32'd33199: dataIn1 = 32'd26
; 
32'd33200: dataIn1 = 32'd27
; 
32'd33201: dataIn1 = 32'd28
; 
32'd33202: dataIn1 = 32'd29
; 
32'd33203: dataIn1 = 32'd30
; 
32'd33204: dataIn1 = 32'd31
; 
32'd33205: dataIn1 = 32'd32
; 
32'd33206: dataIn1 = 32'd33
; 
32'd33207: dataIn1 = 32'd34
; 
32'd33208: dataIn1 = 32'd35
; 
32'd33209: dataIn1 = 32'd36
; 
32'd33210: dataIn1 = 32'd37
; 
32'd33211: dataIn1 = 32'd38
; 
32'd33212: dataIn1 = 32'd40
; 
32'd33213: dataIn1 = 32'd44
; 
32'd33214: dataIn1 = 32'd45
; 
32'd33215: dataIn1 = 32'd46
; 
32'd33216: dataIn1 = 32'd49
; 
32'd33217: dataIn1 = 32'd52
; 
32'd33218: dataIn1 = 32'd53
; 
32'd33219: dataIn1 = 32'd54
; 
32'd33220: dataIn1 = 32'd55
; 
32'd33221: dataIn1 = 32'd56
; 
32'd33222: dataIn1 = 32'd57
; 
32'd33223: dataIn1 = 32'd58
; 
32'd33224: dataIn1 = 32'd59
; 
32'd33225: dataIn1 = 32'd60
; 
32'd33226: dataIn1 = 32'd62
; 
32'd33227: dataIn1 = 32'd63
; 
32'd33228: dataIn1 = 32'd1
; 
32'd33229: dataIn1 = 32'd2
; 
32'd33230: dataIn1 = 32'd3
; 
32'd33231: dataIn1 = 32'd4
; 
32'd33232: dataIn1 = 32'd7
; 
32'd33233: dataIn1 = 32'd8
; 
32'd33234: dataIn1 = 32'd11
; 
32'd33235: dataIn1 = 32'd12
; 
32'd33236: dataIn1 = 32'd14
; 
32'd33237: dataIn1 = 32'd16
; 
32'd33238: dataIn1 = 32'd17
; 
32'd33239: dataIn1 = 32'd18
; 
32'd33240: dataIn1 = 32'd20
; 
32'd33241: dataIn1 = 32'd21
; 
32'd33242: dataIn1 = 32'd22
; 
32'd33243: dataIn1 = 32'd23
; 
32'd33244: dataIn1 = 32'd24
; 
32'd33245: dataIn1 = 32'd26
; 
32'd33246: dataIn1 = 32'd28
; 
32'd33247: dataIn1 = 32'd30
; 
32'd33248: dataIn1 = 32'd31
; 
32'd33249: dataIn1 = 32'd32
; 
32'd33250: dataIn1 = 32'd33
; 
32'd33251: dataIn1 = 32'd34
; 
32'd33252: dataIn1 = 32'd37
; 
32'd33253: dataIn1 = 32'd40
; 
32'd33254: dataIn1 = 32'd41
; 
32'd33255: dataIn1 = 32'd42
; 
32'd33256: dataIn1 = 32'd44
; 
32'd33257: dataIn1 = 32'd46
; 
32'd33258: dataIn1 = 32'd48
; 
32'd33259: dataIn1 = 32'd50
; 
32'd33260: dataIn1 = 32'd51
; 
32'd33261: dataIn1 = 32'd52
; 
32'd33262: dataIn1 = 32'd53
; 
32'd33263: dataIn1 = 32'd54
; 
32'd33264: dataIn1 = 32'd56
; 
32'd33265: dataIn1 = 32'd57
; 
32'd33266: dataIn1 = 32'd60
; 
32'd33267: dataIn1 = 32'd61
; 
32'd33268: dataIn1 = 32'd63
; 
32'd33269: dataIn1 = 32'd0
; 
32'd33270: dataIn1 = 32'd2
; 
32'd33271: dataIn1 = 32'd3
; 
32'd33272: dataIn1 = 32'd4
; 
32'd33273: dataIn1 = 32'd5
; 
32'd33274: dataIn1 = 32'd7
; 
32'd33275: dataIn1 = 32'd10
; 
32'd33276: dataIn1 = 32'd11
; 
32'd33277: dataIn1 = 32'd12
; 
32'd33278: dataIn1 = 32'd13
; 
32'd33279: dataIn1 = 32'd14
; 
32'd33280: dataIn1 = 32'd15
; 
32'd33281: dataIn1 = 32'd16
; 
32'd33282: dataIn1 = 32'd17
; 
32'd33283: dataIn1 = 32'd18
; 
32'd33284: dataIn1 = 32'd19
; 
32'd33285: dataIn1 = 32'd20
; 
32'd33286: dataIn1 = 32'd22
; 
32'd33287: dataIn1 = 32'd24
; 
32'd33288: dataIn1 = 32'd25
; 
32'd33289: dataIn1 = 32'd26
; 
32'd33290: dataIn1 = 32'd29
; 
32'd33291: dataIn1 = 32'd31
; 
32'd33292: dataIn1 = 32'd32
; 
32'd33293: dataIn1 = 32'd33
; 
32'd33294: dataIn1 = 32'd34
; 
32'd33295: dataIn1 = 32'd35
; 
32'd33296: dataIn1 = 32'd39
; 
32'd33297: dataIn1 = 32'd40
; 
32'd33298: dataIn1 = 32'd41
; 
32'd33299: dataIn1 = 32'd42
; 
32'd33300: dataIn1 = 32'd44
; 
32'd33301: dataIn1 = 32'd46
; 
32'd33302: dataIn1 = 32'd47
; 
32'd33303: dataIn1 = 32'd48
; 
32'd33304: dataIn1 = 32'd49
; 
32'd33305: dataIn1 = 32'd51
; 
32'd33306: dataIn1 = 32'd52
; 
32'd33307: dataIn1 = 32'd53
; 
32'd33308: dataIn1 = 32'd55
; 
32'd33309: dataIn1 = 32'd56
; 
32'd33310: dataIn1 = 32'd57
; 
32'd33311: dataIn1 = 32'd58
; 
32'd33312: dataIn1 = 32'd59
; 
32'd33313: dataIn1 = 32'd60
; 
32'd33314: dataIn1 = 32'd61
; 
32'd33315: dataIn1 = 32'd62
; 
32'd33316: dataIn1 = 32'd63
; 
32'd33317: dataIn1 = 32'd0
; 
32'd33318: dataIn1 = 32'd2
; 
32'd33319: dataIn1 = 32'd3
; 
32'd33320: dataIn1 = 32'd4
; 
32'd33321: dataIn1 = 32'd5
; 
32'd33322: dataIn1 = 32'd6
; 
32'd33323: dataIn1 = 32'd7
; 
32'd33324: dataIn1 = 32'd8
; 
32'd33325: dataIn1 = 32'd9
; 
32'd33326: dataIn1 = 32'd10
; 
32'd33327: dataIn1 = 32'd12
; 
32'd33328: dataIn1 = 32'd14
; 
32'd33329: dataIn1 = 32'd17
; 
32'd33330: dataIn1 = 32'd18
; 
32'd33331: dataIn1 = 32'd19
; 
32'd33332: dataIn1 = 32'd22
; 
32'd33333: dataIn1 = 32'd23
; 
32'd33334: dataIn1 = 32'd24
; 
32'd33335: dataIn1 = 32'd26
; 
32'd33336: dataIn1 = 32'd27
; 
32'd33337: dataIn1 = 32'd28
; 
32'd33338: dataIn1 = 32'd29
; 
32'd33339: dataIn1 = 32'd30
; 
32'd33340: dataIn1 = 32'd35
; 
32'd33341: dataIn1 = 32'd36
; 
32'd33342: dataIn1 = 32'd39
; 
32'd33343: dataIn1 = 32'd40
; 
32'd33344: dataIn1 = 32'd41
; 
32'd33345: dataIn1 = 32'd42
; 
32'd33346: dataIn1 = 32'd43
; 
32'd33347: dataIn1 = 32'd44
; 
32'd33348: dataIn1 = 32'd45
; 
32'd33349: dataIn1 = 32'd46
; 
32'd33350: dataIn1 = 32'd47
; 
32'd33351: dataIn1 = 32'd49
; 
32'd33352: dataIn1 = 32'd52
; 
32'd33353: dataIn1 = 32'd53
; 
32'd33354: dataIn1 = 32'd55
; 
32'd33355: dataIn1 = 32'd56
; 
32'd33356: dataIn1 = 32'd57
; 
32'd33357: dataIn1 = 32'd58
; 
32'd33358: dataIn1 = 32'd59
; 
32'd33359: dataIn1 = 32'd61
; 
32'd33360: dataIn1 = 32'd62
; 
32'd33361: dataIn1 = 32'd63
; 
32'd33362: dataIn1 = 32'd0
; 
32'd33363: dataIn1 = 32'd2
; 
32'd33364: dataIn1 = 32'd4
; 
32'd33365: dataIn1 = 32'd5
; 
32'd33366: dataIn1 = 32'd6
; 
32'd33367: dataIn1 = 32'd7
; 
32'd33368: dataIn1 = 32'd9
; 
32'd33369: dataIn1 = 32'd10
; 
32'd33370: dataIn1 = 32'd11
; 
32'd33371: dataIn1 = 32'd14
; 
32'd33372: dataIn1 = 32'd15
; 
32'd33373: dataIn1 = 32'd17
; 
32'd33374: dataIn1 = 32'd18
; 
32'd33375: dataIn1 = 32'd19
; 
32'd33376: dataIn1 = 32'd21
; 
32'd33377: dataIn1 = 32'd22
; 
32'd33378: dataIn1 = 32'd23
; 
32'd33379: dataIn1 = 32'd24
; 
32'd33380: dataIn1 = 32'd25
; 
32'd33381: dataIn1 = 32'd26
; 
32'd33382: dataIn1 = 32'd27
; 
32'd33383: dataIn1 = 32'd28
; 
32'd33384: dataIn1 = 32'd30
; 
32'd33385: dataIn1 = 32'd33
; 
32'd33386: dataIn1 = 32'd35
; 
32'd33387: dataIn1 = 32'd38
; 
32'd33388: dataIn1 = 32'd39
; 
32'd33389: dataIn1 = 32'd42
; 
32'd33390: dataIn1 = 32'd44
; 
32'd33391: dataIn1 = 32'd45
; 
32'd33392: dataIn1 = 32'd46
; 
32'd33393: dataIn1 = 32'd47
; 
32'd33394: dataIn1 = 32'd48
; 
32'd33395: dataIn1 = 32'd49
; 
32'd33396: dataIn1 = 32'd51
; 
32'd33397: dataIn1 = 32'd52
; 
32'd33398: dataIn1 = 32'd53
; 
32'd33399: dataIn1 = 32'd54
; 
32'd33400: dataIn1 = 32'd55
; 
32'd33401: dataIn1 = 32'd56
; 
32'd33402: dataIn1 = 32'd57
; 
32'd33403: dataIn1 = 32'd58
; 
32'd33404: dataIn1 = 32'd59
; 
32'd33405: dataIn1 = 32'd63
; 
32'd33406: dataIn1 = 32'd0
; 
32'd33407: dataIn1 = 32'd1
; 
32'd33408: dataIn1 = 32'd2
; 
32'd33409: dataIn1 = 32'd3
; 
32'd33410: dataIn1 = 32'd5
; 
32'd33411: dataIn1 = 32'd6
; 
32'd33412: dataIn1 = 32'd9
; 
32'd33413: dataIn1 = 32'd10
; 
32'd33414: dataIn1 = 32'd11
; 
32'd33415: dataIn1 = 32'd12
; 
32'd33416: dataIn1 = 32'd13
; 
32'd33417: dataIn1 = 32'd16
; 
32'd33418: dataIn1 = 32'd17
; 
32'd33419: dataIn1 = 32'd18
; 
32'd33420: dataIn1 = 32'd19
; 
32'd33421: dataIn1 = 32'd20
; 
32'd33422: dataIn1 = 32'd21
; 
32'd33423: dataIn1 = 32'd22
; 
32'd33424: dataIn1 = 32'd24
; 
32'd33425: dataIn1 = 32'd25
; 
32'd33426: dataIn1 = 32'd26
; 
32'd33427: dataIn1 = 32'd27
; 
32'd33428: dataIn1 = 32'd28
; 
32'd33429: dataIn1 = 32'd29
; 
32'd33430: dataIn1 = 32'd32
; 
32'd33431: dataIn1 = 32'd33
; 
32'd33432: dataIn1 = 32'd35
; 
32'd33433: dataIn1 = 32'd36
; 
32'd33434: dataIn1 = 32'd37
; 
32'd33435: dataIn1 = 32'd39
; 
32'd33436: dataIn1 = 32'd41
; 
32'd33437: dataIn1 = 32'd43
; 
32'd33438: dataIn1 = 32'd44
; 
32'd33439: dataIn1 = 32'd45
; 
32'd33440: dataIn1 = 32'd46
; 
32'd33441: dataIn1 = 32'd47
; 
32'd33442: dataIn1 = 32'd49
; 
32'd33443: dataIn1 = 32'd56
; 
32'd33444: dataIn1 = 32'd57
; 
32'd33445: dataIn1 = 32'd59
; 
32'd33446: dataIn1 = 32'd61
; 
32'd33447: dataIn1 = 32'd62
; 
32'd33448: dataIn1 = 32'd0
; 
32'd33449: dataIn1 = 32'd1
; 
32'd33450: dataIn1 = 32'd2
; 
32'd33451: dataIn1 = 32'd6
; 
32'd33452: dataIn1 = 32'd7
; 
32'd33453: dataIn1 = 32'd11
; 
32'd33454: dataIn1 = 32'd13
; 
32'd33455: dataIn1 = 32'd14
; 
32'd33456: dataIn1 = 32'd20
; 
32'd33457: dataIn1 = 32'd21
; 
32'd33458: dataIn1 = 32'd26
; 
32'd33459: dataIn1 = 32'd27
; 
32'd33460: dataIn1 = 32'd28
; 
32'd33461: dataIn1 = 32'd31
; 
32'd33462: dataIn1 = 32'd32
; 
32'd33463: dataIn1 = 32'd33
; 
32'd33464: dataIn1 = 32'd35
; 
32'd33465: dataIn1 = 32'd37
; 
32'd33466: dataIn1 = 32'd38
; 
32'd33467: dataIn1 = 32'd39
; 
32'd33468: dataIn1 = 32'd42
; 
32'd33469: dataIn1 = 32'd45
; 
32'd33470: dataIn1 = 32'd47
; 
32'd33471: dataIn1 = 32'd48
; 
32'd33472: dataIn1 = 32'd50
; 
32'd33473: dataIn1 = 32'd51
; 
32'd33474: dataIn1 = 32'd52
; 
32'd33475: dataIn1 = 32'd55
; 
32'd33476: dataIn1 = 32'd56
; 
32'd33477: dataIn1 = 32'd57
; 
32'd33478: dataIn1 = 32'd58
; 
32'd33479: dataIn1 = 32'd59
; 
32'd33480: dataIn1 = 32'd60
; 
32'd33481: dataIn1 = 32'd62
; 
32'd33482: dataIn1 = 32'd63
; 
32'd33483: dataIn1 = 32'd0
; 
32'd33484: dataIn1 = 32'd2
; 
32'd33485: dataIn1 = 32'd3
; 
32'd33486: dataIn1 = 32'd6
; 
32'd33487: dataIn1 = 32'd7
; 
32'd33488: dataIn1 = 32'd8
; 
32'd33489: dataIn1 = 32'd10
; 
32'd33490: dataIn1 = 32'd11
; 
32'd33491: dataIn1 = 32'd12
; 
32'd33492: dataIn1 = 32'd14
; 
32'd33493: dataIn1 = 32'd17
; 
32'd33494: dataIn1 = 32'd19
; 
32'd33495: dataIn1 = 32'd20
; 
32'd33496: dataIn1 = 32'd21
; 
32'd33497: dataIn1 = 32'd22
; 
32'd33498: dataIn1 = 32'd23
; 
32'd33499: dataIn1 = 32'd24
; 
32'd33500: dataIn1 = 32'd25
; 
32'd33501: dataIn1 = 32'd26
; 
32'd33502: dataIn1 = 32'd29
; 
32'd33503: dataIn1 = 32'd30
; 
32'd33504: dataIn1 = 32'd33
; 
32'd33505: dataIn1 = 32'd34
; 
32'd33506: dataIn1 = 32'd35
; 
32'd33507: dataIn1 = 32'd36
; 
32'd33508: dataIn1 = 32'd37
; 
32'd33509: dataIn1 = 32'd38
; 
32'd33510: dataIn1 = 32'd39
; 
32'd33511: dataIn1 = 32'd40
; 
32'd33512: dataIn1 = 32'd41
; 
32'd33513: dataIn1 = 32'd42
; 
32'd33514: dataIn1 = 32'd44
; 
32'd33515: dataIn1 = 32'd46
; 
32'd33516: dataIn1 = 32'd47
; 
32'd33517: dataIn1 = 32'd49
; 
32'd33518: dataIn1 = 32'd50
; 
32'd33519: dataIn1 = 32'd51
; 
32'd33520: dataIn1 = 32'd53
; 
32'd33521: dataIn1 = 32'd56
; 
32'd33522: dataIn1 = 32'd58
; 
32'd33523: dataIn1 = 32'd59
; 
32'd33524: dataIn1 = 32'd61
; 
32'd33525: dataIn1 = 32'd62
; 
32'd33526: dataIn1 = 32'd63
; 
32'd33527: dataIn1 = 32'd1
; 
32'd33528: dataIn1 = 32'd2
; 
32'd33529: dataIn1 = 32'd3
; 
32'd33530: dataIn1 = 32'd4
; 
32'd33531: dataIn1 = 32'd5
; 
32'd33532: dataIn1 = 32'd12
; 
32'd33533: dataIn1 = 32'd14
; 
32'd33534: dataIn1 = 32'd15
; 
32'd33535: dataIn1 = 32'd16
; 
32'd33536: dataIn1 = 32'd19
; 
32'd33537: dataIn1 = 32'd20
; 
32'd33538: dataIn1 = 32'd21
; 
32'd33539: dataIn1 = 32'd22
; 
32'd33540: dataIn1 = 32'd23
; 
32'd33541: dataIn1 = 32'd24
; 
32'd33542: dataIn1 = 32'd25
; 
32'd33543: dataIn1 = 32'd26
; 
32'd33544: dataIn1 = 32'd28
; 
32'd33545: dataIn1 = 32'd29
; 
32'd33546: dataIn1 = 32'd30
; 
32'd33547: dataIn1 = 32'd33
; 
32'd33548: dataIn1 = 32'd34
; 
32'd33549: dataIn1 = 32'd35
; 
32'd33550: dataIn1 = 32'd37
; 
32'd33551: dataIn1 = 32'd39
; 
32'd33552: dataIn1 = 32'd40
; 
32'd33553: dataIn1 = 32'd43
; 
32'd33554: dataIn1 = 32'd45
; 
32'd33555: dataIn1 = 32'd49
; 
32'd33556: dataIn1 = 32'd50
; 
32'd33557: dataIn1 = 32'd52
; 
32'd33558: dataIn1 = 32'd53
; 
32'd33559: dataIn1 = 32'd54
; 
32'd33560: dataIn1 = 32'd55
; 
32'd33561: dataIn1 = 32'd56
; 
32'd33562: dataIn1 = 32'd57
; 
32'd33563: dataIn1 = 32'd58
; 
32'd33564: dataIn1 = 32'd59
; 
32'd33565: dataIn1 = 32'd60
; 
32'd33566: dataIn1 = 32'd61
; 
32'd33567: dataIn1 = 32'd62
; 
32'd33568: dataIn1 = 32'd63
; 
32'd33569: dataIn1 = 32'd0
; 
32'd33570: dataIn1 = 32'd1
; 
32'd33571: dataIn1 = 32'd3
; 
32'd33572: dataIn1 = 32'd4
; 
32'd33573: dataIn1 = 32'd6
; 
32'd33574: dataIn1 = 32'd7
; 
32'd33575: dataIn1 = 32'd8
; 
32'd33576: dataIn1 = 32'd10
; 
32'd33577: dataIn1 = 32'd11
; 
32'd33578: dataIn1 = 32'd12
; 
32'd33579: dataIn1 = 32'd13
; 
32'd33580: dataIn1 = 32'd14
; 
32'd33581: dataIn1 = 32'd15
; 
32'd33582: dataIn1 = 32'd19
; 
32'd33583: dataIn1 = 32'd20
; 
32'd33584: dataIn1 = 32'd21
; 
32'd33585: dataIn1 = 32'd22
; 
32'd33586: dataIn1 = 32'd23
; 
32'd33587: dataIn1 = 32'd24
; 
32'd33588: dataIn1 = 32'd25
; 
32'd33589: dataIn1 = 32'd26
; 
32'd33590: dataIn1 = 32'd29
; 
32'd33591: dataIn1 = 32'd31
; 
32'd33592: dataIn1 = 32'd33
; 
32'd33593: dataIn1 = 32'd34
; 
32'd33594: dataIn1 = 32'd35
; 
32'd33595: dataIn1 = 32'd36
; 
32'd33596: dataIn1 = 32'd37
; 
32'd33597: dataIn1 = 32'd38
; 
32'd33598: dataIn1 = 32'd39
; 
32'd33599: dataIn1 = 32'd41
; 
32'd33600: dataIn1 = 32'd43
; 
32'd33601: dataIn1 = 32'd44
; 
32'd33602: dataIn1 = 32'd46
; 
32'd33603: dataIn1 = 32'd47
; 
32'd33604: dataIn1 = 32'd48
; 
32'd33605: dataIn1 = 32'd49
; 
32'd33606: dataIn1 = 32'd51
; 
32'd33607: dataIn1 = 32'd52
; 
32'd33608: dataIn1 = 32'd56
; 
32'd33609: dataIn1 = 32'd57
; 
32'd33610: dataIn1 = 32'd59
; 
32'd33611: dataIn1 = 32'd60
; 
32'd33612: dataIn1 = 32'd62
; 
32'd33613: dataIn1 = 32'd0
; 
32'd33614: dataIn1 = 32'd2
; 
32'd33615: dataIn1 = 32'd3
; 
32'd33616: dataIn1 = 32'd4
; 
32'd33617: dataIn1 = 32'd6
; 
32'd33618: dataIn1 = 32'd7
; 
32'd33619: dataIn1 = 32'd8
; 
32'd33620: dataIn1 = 32'd9
; 
32'd33621: dataIn1 = 32'd10
; 
32'd33622: dataIn1 = 32'd13
; 
32'd33623: dataIn1 = 32'd16
; 
32'd33624: dataIn1 = 32'd17
; 
32'd33625: dataIn1 = 32'd18
; 
32'd33626: dataIn1 = 32'd19
; 
32'd33627: dataIn1 = 32'd20
; 
32'd33628: dataIn1 = 32'd21
; 
32'd33629: dataIn1 = 32'd22
; 
32'd33630: dataIn1 = 32'd23
; 
32'd33631: dataIn1 = 32'd24
; 
32'd33632: dataIn1 = 32'd27
; 
32'd33633: dataIn1 = 32'd28
; 
32'd33634: dataIn1 = 32'd29
; 
32'd33635: dataIn1 = 32'd31
; 
32'd33636: dataIn1 = 32'd32
; 
32'd33637: dataIn1 = 32'd34
; 
32'd33638: dataIn1 = 32'd35
; 
32'd33639: dataIn1 = 32'd36
; 
32'd33640: dataIn1 = 32'd37
; 
32'd33641: dataIn1 = 32'd40
; 
32'd33642: dataIn1 = 32'd41
; 
32'd33643: dataIn1 = 32'd42
; 
32'd33644: dataIn1 = 32'd43
; 
32'd33645: dataIn1 = 32'd44
; 
32'd33646: dataIn1 = 32'd45
; 
32'd33647: dataIn1 = 32'd47
; 
32'd33648: dataIn1 = 32'd48
; 
32'd33649: dataIn1 = 32'd49
; 
32'd33650: dataIn1 = 32'd50
; 
32'd33651: dataIn1 = 32'd51
; 
32'd33652: dataIn1 = 32'd53
; 
32'd33653: dataIn1 = 32'd54
; 
32'd33654: dataIn1 = 32'd55
; 
32'd33655: dataIn1 = 32'd56
; 
32'd33656: dataIn1 = 32'd58
; 
32'd33657: dataIn1 = 32'd59
; 
32'd33658: dataIn1 = 32'd61
; 
32'd33659: dataIn1 = 32'd1
; 
32'd33660: dataIn1 = 32'd2
; 
32'd33661: dataIn1 = 32'd3
; 
32'd33662: dataIn1 = 32'd4
; 
32'd33663: dataIn1 = 32'd5
; 
32'd33664: dataIn1 = 32'd6
; 
32'd33665: dataIn1 = 32'd7
; 
32'd33666: dataIn1 = 32'd8
; 
32'd33667: dataIn1 = 32'd9
; 
32'd33668: dataIn1 = 32'd11
; 
32'd33669: dataIn1 = 32'd12
; 
32'd33670: dataIn1 = 32'd13
; 
32'd33671: dataIn1 = 32'd14
; 
32'd33672: dataIn1 = 32'd17
; 
32'd33673: dataIn1 = 32'd18
; 
32'd33674: dataIn1 = 32'd19
; 
32'd33675: dataIn1 = 32'd20
; 
32'd33676: dataIn1 = 32'd21
; 
32'd33677: dataIn1 = 32'd26
; 
32'd33678: dataIn1 = 32'd27
; 
32'd33679: dataIn1 = 32'd28
; 
32'd33680: dataIn1 = 32'd29
; 
32'd33681: dataIn1 = 32'd31
; 
32'd33682: dataIn1 = 32'd32
; 
32'd33683: dataIn1 = 32'd33
; 
32'd33684: dataIn1 = 32'd36
; 
32'd33685: dataIn1 = 32'd38
; 
32'd33686: dataIn1 = 32'd39
; 
32'd33687: dataIn1 = 32'd40
; 
32'd33688: dataIn1 = 32'd42
; 
32'd33689: dataIn1 = 32'd43
; 
32'd33690: dataIn1 = 32'd45
; 
32'd33691: dataIn1 = 32'd46
; 
32'd33692: dataIn1 = 32'd47
; 
32'd33693: dataIn1 = 32'd48
; 
32'd33694: dataIn1 = 32'd50
; 
32'd33695: dataIn1 = 32'd51
; 
32'd33696: dataIn1 = 32'd54
; 
32'd33697: dataIn1 = 32'd55
; 
32'd33698: dataIn1 = 32'd57
; 
32'd33699: dataIn1 = 32'd59
; 
32'd33700: dataIn1 = 32'd61
; 
32'd33701: dataIn1 = 32'd62
; 
32'd33702: dataIn1 = 32'd63
; 
32'd33703: dataIn1 = 32'd0
; 
32'd33704: dataIn1 = 32'd1
; 
32'd33705: dataIn1 = 32'd4
; 
32'd33706: dataIn1 = 32'd5
; 
32'd33707: dataIn1 = 32'd6
; 
32'd33708: dataIn1 = 32'd8
; 
32'd33709: dataIn1 = 32'd9
; 
32'd33710: dataIn1 = 32'd10
; 
32'd33711: dataIn1 = 32'd11
; 
32'd33712: dataIn1 = 32'd14
; 
32'd33713: dataIn1 = 32'd21
; 
32'd33714: dataIn1 = 32'd22
; 
32'd33715: dataIn1 = 32'd23
; 
32'd33716: dataIn1 = 32'd26
; 
32'd33717: dataIn1 = 32'd27
; 
32'd33718: dataIn1 = 32'd29
; 
32'd33719: dataIn1 = 32'd30
; 
32'd33720: dataIn1 = 32'd31
; 
32'd33721: dataIn1 = 32'd33
; 
32'd33722: dataIn1 = 32'd34
; 
32'd33723: dataIn1 = 32'd35
; 
32'd33724: dataIn1 = 32'd37
; 
32'd33725: dataIn1 = 32'd38
; 
32'd33726: dataIn1 = 32'd39
; 
32'd33727: dataIn1 = 32'd40
; 
32'd33728: dataIn1 = 32'd41
; 
32'd33729: dataIn1 = 32'd42
; 
32'd33730: dataIn1 = 32'd43
; 
32'd33731: dataIn1 = 32'd44
; 
32'd33732: dataIn1 = 32'd46
; 
32'd33733: dataIn1 = 32'd47
; 
32'd33734: dataIn1 = 32'd48
; 
32'd33735: dataIn1 = 32'd50
; 
32'd33736: dataIn1 = 32'd51
; 
32'd33737: dataIn1 = 32'd52
; 
32'd33738: dataIn1 = 32'd55
; 
32'd33739: dataIn1 = 32'd56
; 
32'd33740: dataIn1 = 32'd57
; 
32'd33741: dataIn1 = 32'd59
; 
32'd33742: dataIn1 = 32'd60
; 
32'd33743: dataIn1 = 32'd62
; 
32'd33744: dataIn1 = 32'd0
; 
32'd33745: dataIn1 = 32'd1
; 
32'd33746: dataIn1 = 32'd2
; 
32'd33747: dataIn1 = 32'd4
; 
32'd33748: dataIn1 = 32'd6
; 
32'd33749: dataIn1 = 32'd7
; 
32'd33750: dataIn1 = 32'd10
; 
32'd33751: dataIn1 = 32'd12
; 
32'd33752: dataIn1 = 32'd13
; 
32'd33753: dataIn1 = 32'd14
; 
32'd33754: dataIn1 = 32'd15
; 
32'd33755: dataIn1 = 32'd17
; 
32'd33756: dataIn1 = 32'd18
; 
32'd33757: dataIn1 = 32'd19
; 
32'd33758: dataIn1 = 32'd20
; 
32'd33759: dataIn1 = 32'd22
; 
32'd33760: dataIn1 = 32'd23
; 
32'd33761: dataIn1 = 32'd26
; 
32'd33762: dataIn1 = 32'd27
; 
32'd33763: dataIn1 = 32'd28
; 
32'd33764: dataIn1 = 32'd29
; 
32'd33765: dataIn1 = 32'd30
; 
32'd33766: dataIn1 = 32'd31
; 
32'd33767: dataIn1 = 32'd33
; 
32'd33768: dataIn1 = 32'd34
; 
32'd33769: dataIn1 = 32'd36
; 
32'd33770: dataIn1 = 32'd40
; 
32'd33771: dataIn1 = 32'd42
; 
32'd33772: dataIn1 = 32'd43
; 
32'd33773: dataIn1 = 32'd47
; 
32'd33774: dataIn1 = 32'd48
; 
32'd33775: dataIn1 = 32'd49
; 
32'd33776: dataIn1 = 32'd50
; 
32'd33777: dataIn1 = 32'd51
; 
32'd33778: dataIn1 = 32'd52
; 
32'd33779: dataIn1 = 32'd55
; 
32'd33780: dataIn1 = 32'd56
; 
32'd33781: dataIn1 = 32'd57
; 
32'd33782: dataIn1 = 32'd58
; 
32'd33783: dataIn1 = 32'd59
; 
32'd33784: dataIn1 = 32'd60
; 
32'd33785: dataIn1 = 32'd61
; 
32'd33786: dataIn1 = 32'd62
; 
32'd33787: dataIn1 = 32'd63
; 
32'd33788: dataIn1 = 32'd2
; 
32'd33789: dataIn1 = 32'd3
; 
32'd33790: dataIn1 = 32'd5
; 
32'd33791: dataIn1 = 32'd7
; 
32'd33792: dataIn1 = 32'd9
; 
32'd33793: dataIn1 = 32'd10
; 
32'd33794: dataIn1 = 32'd12
; 
32'd33795: dataIn1 = 32'd13
; 
32'd33796: dataIn1 = 32'd18
; 
32'd33797: dataIn1 = 32'd19
; 
32'd33798: dataIn1 = 32'd20
; 
32'd33799: dataIn1 = 32'd21
; 
32'd33800: dataIn1 = 32'd22
; 
32'd33801: dataIn1 = 32'd23
; 
32'd33802: dataIn1 = 32'd24
; 
32'd33803: dataIn1 = 32'd26
; 
32'd33804: dataIn1 = 32'd27
; 
32'd33805: dataIn1 = 32'd28
; 
32'd33806: dataIn1 = 32'd29
; 
32'd33807: dataIn1 = 32'd30
; 
32'd33808: dataIn1 = 32'd32
; 
32'd33809: dataIn1 = 32'd34
; 
32'd33810: dataIn1 = 32'd35
; 
32'd33811: dataIn1 = 32'd37
; 
32'd33812: dataIn1 = 32'd38
; 
32'd33813: dataIn1 = 32'd39
; 
32'd33814: dataIn1 = 32'd40
; 
32'd33815: dataIn1 = 32'd41
; 
32'd33816: dataIn1 = 32'd43
; 
32'd33817: dataIn1 = 32'd44
; 
32'd33818: dataIn1 = 32'd45
; 
32'd33819: dataIn1 = 32'd47
; 
32'd33820: dataIn1 = 32'd49
; 
32'd33821: dataIn1 = 32'd50
; 
32'd33822: dataIn1 = 32'd51
; 
32'd33823: dataIn1 = 32'd52
; 
32'd33824: dataIn1 = 32'd53
; 
32'd33825: dataIn1 = 32'd55
; 
32'd33826: dataIn1 = 32'd56
; 
32'd33827: dataIn1 = 32'd57
; 
32'd33828: dataIn1 = 32'd59
; 
32'd33829: dataIn1 = 32'd60
; 
32'd33830: dataIn1 = 32'd61
; 
32'd33831: dataIn1 = 32'd62
; 
32'd33832: dataIn1 = 32'd0
; 
32'd33833: dataIn1 = 32'd1
; 
32'd33834: dataIn1 = 32'd2
; 
32'd33835: dataIn1 = 32'd3
; 
32'd33836: dataIn1 = 32'd4
; 
32'd33837: dataIn1 = 32'd5
; 
32'd33838: dataIn1 = 32'd7
; 
32'd33839: dataIn1 = 32'd9
; 
32'd33840: dataIn1 = 32'd11
; 
32'd33841: dataIn1 = 32'd12
; 
32'd33842: dataIn1 = 32'd13
; 
32'd33843: dataIn1 = 32'd14
; 
32'd33844: dataIn1 = 32'd15
; 
32'd33845: dataIn1 = 32'd16
; 
32'd33846: dataIn1 = 32'd17
; 
32'd33847: dataIn1 = 32'd18
; 
32'd33848: dataIn1 = 32'd19
; 
32'd33849: dataIn1 = 32'd20
; 
32'd33850: dataIn1 = 32'd21
; 
32'd33851: dataIn1 = 32'd22
; 
32'd33852: dataIn1 = 32'd23
; 
32'd33853: dataIn1 = 32'd24
; 
32'd33854: dataIn1 = 32'd25
; 
32'd33855: dataIn1 = 32'd26
; 
32'd33856: dataIn1 = 32'd28
; 
32'd33857: dataIn1 = 32'd29
; 
32'd33858: dataIn1 = 32'd30
; 
32'd33859: dataIn1 = 32'd31
; 
32'd33860: dataIn1 = 32'd32
; 
32'd33861: dataIn1 = 32'd33
; 
32'd33862: dataIn1 = 32'd40
; 
32'd33863: dataIn1 = 32'd41
; 
32'd33864: dataIn1 = 32'd43
; 
32'd33865: dataIn1 = 32'd44
; 
32'd33866: dataIn1 = 32'd45
; 
32'd33867: dataIn1 = 32'd46
; 
32'd33868: dataIn1 = 32'd47
; 
32'd33869: dataIn1 = 32'd49
; 
32'd33870: dataIn1 = 32'd52
; 
32'd33871: dataIn1 = 32'd57
; 
32'd33872: dataIn1 = 32'd59
; 
32'd33873: dataIn1 = 32'd60
; 
32'd33874: dataIn1 = 32'd61
; 
32'd33875: dataIn1 = 32'd62
; 
32'd33876: dataIn1 = 32'd3
; 
32'd33877: dataIn1 = 32'd4
; 
32'd33878: dataIn1 = 32'd5
; 
32'd33879: dataIn1 = 32'd6
; 
32'd33880: dataIn1 = 32'd10
; 
32'd33881: dataIn1 = 32'd11
; 
32'd33882: dataIn1 = 32'd12
; 
32'd33883: dataIn1 = 32'd13
; 
32'd33884: dataIn1 = 32'd14
; 
32'd33885: dataIn1 = 32'd15
; 
32'd33886: dataIn1 = 32'd16
; 
32'd33887: dataIn1 = 32'd18
; 
32'd33888: dataIn1 = 32'd20
; 
32'd33889: dataIn1 = 32'd21
; 
32'd33890: dataIn1 = 32'd22
; 
32'd33891: dataIn1 = 32'd23
; 
32'd33892: dataIn1 = 32'd24
; 
32'd33893: dataIn1 = 32'd25
; 
32'd33894: dataIn1 = 32'd27
; 
32'd33895: dataIn1 = 32'd28
; 
32'd33896: dataIn1 = 32'd29
; 
32'd33897: dataIn1 = 32'd31
; 
32'd33898: dataIn1 = 32'd32
; 
32'd33899: dataIn1 = 32'd33
; 
32'd33900: dataIn1 = 32'd34
; 
32'd33901: dataIn1 = 32'd36
; 
32'd33902: dataIn1 = 32'd37
; 
32'd33903: dataIn1 = 32'd38
; 
32'd33904: dataIn1 = 32'd40
; 
32'd33905: dataIn1 = 32'd42
; 
32'd33906: dataIn1 = 32'd45
; 
32'd33907: dataIn1 = 32'd46
; 
32'd33908: dataIn1 = 32'd47
; 
32'd33909: dataIn1 = 32'd50
; 
32'd33910: dataIn1 = 32'd51
; 
32'd33911: dataIn1 = 32'd52
; 
32'd33912: dataIn1 = 32'd53
; 
32'd33913: dataIn1 = 32'd54
; 
32'd33914: dataIn1 = 32'd55
; 
32'd33915: dataIn1 = 32'd57
; 
32'd33916: dataIn1 = 32'd58
; 
32'd33917: dataIn1 = 32'd59
; 
32'd33918: dataIn1 = 32'd62
; 
32'd33919: dataIn1 = 32'd63
; 
32'd33920: dataIn1 = 32'd0
; 
32'd33921: dataIn1 = 32'd2
; 
32'd33922: dataIn1 = 32'd3
; 
32'd33923: dataIn1 = 32'd5
; 
32'd33924: dataIn1 = 32'd6
; 
32'd33925: dataIn1 = 32'd8
; 
32'd33926: dataIn1 = 32'd10
; 
32'd33927: dataIn1 = 32'd11
; 
32'd33928: dataIn1 = 32'd14
; 
32'd33929: dataIn1 = 32'd15
; 
32'd33930: dataIn1 = 32'd16
; 
32'd33931: dataIn1 = 32'd17
; 
32'd33932: dataIn1 = 32'd18
; 
32'd33933: dataIn1 = 32'd19
; 
32'd33934: dataIn1 = 32'd21
; 
32'd33935: dataIn1 = 32'd22
; 
32'd33936: dataIn1 = 32'd23
; 
32'd33937: dataIn1 = 32'd25
; 
32'd33938: dataIn1 = 32'd30
; 
32'd33939: dataIn1 = 32'd32
; 
32'd33940: dataIn1 = 32'd33
; 
32'd33941: dataIn1 = 32'd34
; 
32'd33942: dataIn1 = 32'd35
; 
32'd33943: dataIn1 = 32'd36
; 
32'd33944: dataIn1 = 32'd37
; 
32'd33945: dataIn1 = 32'd38
; 
32'd33946: dataIn1 = 32'd39
; 
32'd33947: dataIn1 = 32'd42
; 
32'd33948: dataIn1 = 32'd44
; 
32'd33949: dataIn1 = 32'd46
; 
32'd33950: dataIn1 = 32'd48
; 
32'd33951: dataIn1 = 32'd49
; 
32'd33952: dataIn1 = 32'd50
; 
32'd33953: dataIn1 = 32'd51
; 
32'd33954: dataIn1 = 32'd52
; 
32'd33955: dataIn1 = 32'd55
; 
32'd33956: dataIn1 = 32'd56
; 
32'd33957: dataIn1 = 32'd57
; 
32'd33958: dataIn1 = 32'd58
; 
32'd33959: dataIn1 = 32'd60
; 
32'd33960: dataIn1 = 32'd61
; 
32'd33961: dataIn1 = 32'd62
; 
32'd33962: dataIn1 = 32'd2
; 
32'd33963: dataIn1 = 32'd3
; 
32'd33964: dataIn1 = 32'd4
; 
32'd33965: dataIn1 = 32'd8
; 
32'd33966: dataIn1 = 32'd9
; 
32'd33967: dataIn1 = 32'd10
; 
32'd33968: dataIn1 = 32'd12
; 
32'd33969: dataIn1 = 32'd14
; 
32'd33970: dataIn1 = 32'd17
; 
32'd33971: dataIn1 = 32'd19
; 
32'd33972: dataIn1 = 32'd20
; 
32'd33973: dataIn1 = 32'd21
; 
32'd33974: dataIn1 = 32'd22
; 
32'd33975: dataIn1 = 32'd24
; 
32'd33976: dataIn1 = 32'd27
; 
32'd33977: dataIn1 = 32'd31
; 
32'd33978: dataIn1 = 32'd32
; 
32'd33979: dataIn1 = 32'd33
; 
32'd33980: dataIn1 = 32'd35
; 
32'd33981: dataIn1 = 32'd36
; 
32'd33982: dataIn1 = 32'd38
; 
32'd33983: dataIn1 = 32'd40
; 
32'd33984: dataIn1 = 32'd41
; 
32'd33985: dataIn1 = 32'd42
; 
32'd33986: dataIn1 = 32'd44
; 
32'd33987: dataIn1 = 32'd45
; 
32'd33988: dataIn1 = 32'd46
; 
32'd33989: dataIn1 = 32'd47
; 
32'd33990: dataIn1 = 32'd51
; 
32'd33991: dataIn1 = 32'd53
; 
32'd33992: dataIn1 = 32'd54
; 
32'd33993: dataIn1 = 32'd55
; 
32'd33994: dataIn1 = 32'd56
; 
32'd33995: dataIn1 = 32'd57
; 
32'd33996: dataIn1 = 32'd58
; 
32'd33997: dataIn1 = 32'd60
; 
32'd33998: dataIn1 = 32'd62
; 
32'd33999: dataIn1 = 32'd0
; 
32'd34000: dataIn1 = 32'd3
; 
32'd34001: dataIn1 = 32'd4
; 
32'd34002: dataIn1 = 32'd5
; 
32'd34003: dataIn1 = 32'd6
; 
32'd34004: dataIn1 = 32'd7
; 
32'd34005: dataIn1 = 32'd8
; 
32'd34006: dataIn1 = 32'd9
; 
32'd34007: dataIn1 = 32'd11
; 
32'd34008: dataIn1 = 32'd12
; 
32'd34009: dataIn1 = 32'd13
; 
32'd34010: dataIn1 = 32'd14
; 
32'd34011: dataIn1 = 32'd15
; 
32'd34012: dataIn1 = 32'd17
; 
32'd34013: dataIn1 = 32'd18
; 
32'd34014: dataIn1 = 32'd19
; 
32'd34015: dataIn1 = 32'd21
; 
32'd34016: dataIn1 = 32'd23
; 
32'd34017: dataIn1 = 32'd24
; 
32'd34018: dataIn1 = 32'd25
; 
32'd34019: dataIn1 = 32'd26
; 
32'd34020: dataIn1 = 32'd27
; 
32'd34021: dataIn1 = 32'd29
; 
32'd34022: dataIn1 = 32'd31
; 
32'd34023: dataIn1 = 32'd32
; 
32'd34024: dataIn1 = 32'd34
; 
32'd34025: dataIn1 = 32'd36
; 
32'd34026: dataIn1 = 32'd38
; 
32'd34027: dataIn1 = 32'd40
; 
32'd34028: dataIn1 = 32'd43
; 
32'd34029: dataIn1 = 32'd44
; 
32'd34030: dataIn1 = 32'd45
; 
32'd34031: dataIn1 = 32'd46
; 
32'd34032: dataIn1 = 32'd47
; 
32'd34033: dataIn1 = 32'd48
; 
32'd34034: dataIn1 = 32'd49
; 
32'd34035: dataIn1 = 32'd52
; 
32'd34036: dataIn1 = 32'd53
; 
32'd34037: dataIn1 = 32'd54
; 
32'd34038: dataIn1 = 32'd55
; 
32'd34039: dataIn1 = 32'd56
; 
32'd34040: dataIn1 = 32'd58
; 
32'd34041: dataIn1 = 32'd59
; 
32'd34042: dataIn1 = 32'd60
; 
32'd34043: dataIn1 = 32'd61
; 
32'd34044: dataIn1 = 32'd63
; 
32'd34045: dataIn1 = 32'd0
; 
32'd34046: dataIn1 = 32'd1
; 
32'd34047: dataIn1 = 32'd2
; 
32'd34048: dataIn1 = 32'd5
; 
32'd34049: dataIn1 = 32'd6
; 
32'd34050: dataIn1 = 32'd7
; 
32'd34051: dataIn1 = 32'd8
; 
32'd34052: dataIn1 = 32'd9
; 
32'd34053: dataIn1 = 32'd11
; 
32'd34054: dataIn1 = 32'd14
; 
32'd34055: dataIn1 = 32'd15
; 
32'd34056: dataIn1 = 32'd16
; 
32'd34057: dataIn1 = 32'd17
; 
32'd34058: dataIn1 = 32'd18
; 
32'd34059: dataIn1 = 32'd19
; 
32'd34060: dataIn1 = 32'd20
; 
32'd34061: dataIn1 = 32'd21
; 
32'd34062: dataIn1 = 32'd24
; 
32'd34063: dataIn1 = 32'd25
; 
32'd34064: dataIn1 = 32'd26
; 
32'd34065: dataIn1 = 32'd28
; 
32'd34066: dataIn1 = 32'd30
; 
32'd34067: dataIn1 = 32'd32
; 
32'd34068: dataIn1 = 32'd33
; 
32'd34069: dataIn1 = 32'd36
; 
32'd34070: dataIn1 = 32'd37
; 
32'd34071: dataIn1 = 32'd39
; 
32'd34072: dataIn1 = 32'd41
; 
32'd34073: dataIn1 = 32'd42
; 
32'd34074: dataIn1 = 32'd46
; 
32'd34075: dataIn1 = 32'd47
; 
32'd34076: dataIn1 = 32'd48
; 
32'd34077: dataIn1 = 32'd49
; 
32'd34078: dataIn1 = 32'd50
; 
32'd34079: dataIn1 = 32'd51
; 
32'd34080: dataIn1 = 32'd52
; 
32'd34081: dataIn1 = 32'd55
; 
32'd34082: dataIn1 = 32'd56
; 
32'd34083: dataIn1 = 32'd57
; 
32'd34084: dataIn1 = 32'd58
; 
32'd34085: dataIn1 = 32'd59
; 
32'd34086: dataIn1 = 32'd62
; 
32'd34087: dataIn1 = 32'd63
; 
32'd34088: dataIn1 = 32'd0
; 
32'd34089: dataIn1 = 32'd2
; 
32'd34090: dataIn1 = 32'd3
; 
32'd34091: dataIn1 = 32'd5
; 
32'd34092: dataIn1 = 32'd8
; 
32'd34093: dataIn1 = 32'd9
; 
32'd34094: dataIn1 = 32'd10
; 
32'd34095: dataIn1 = 32'd11
; 
32'd34096: dataIn1 = 32'd12
; 
32'd34097: dataIn1 = 32'd15
; 
32'd34098: dataIn1 = 32'd16
; 
32'd34099: dataIn1 = 32'd17
; 
32'd34100: dataIn1 = 32'd18
; 
32'd34101: dataIn1 = 32'd19
; 
32'd34102: dataIn1 = 32'd21
; 
32'd34103: dataIn1 = 32'd22
; 
32'd34104: dataIn1 = 32'd23
; 
32'd34105: dataIn1 = 32'd24
; 
32'd34106: dataIn1 = 32'd25
; 
32'd34107: dataIn1 = 32'd26
; 
32'd34108: dataIn1 = 32'd27
; 
32'd34109: dataIn1 = 32'd29
; 
32'd34110: dataIn1 = 32'd30
; 
32'd34111: dataIn1 = 32'd31
; 
32'd34112: dataIn1 = 32'd32
; 
32'd34113: dataIn1 = 32'd33
; 
32'd34114: dataIn1 = 32'd35
; 
32'd34115: dataIn1 = 32'd36
; 
32'd34116: dataIn1 = 32'd37
; 
32'd34117: dataIn1 = 32'd40
; 
32'd34118: dataIn1 = 32'd41
; 
32'd34119: dataIn1 = 32'd42
; 
32'd34120: dataIn1 = 32'd43
; 
32'd34121: dataIn1 = 32'd44
; 
32'd34122: dataIn1 = 32'd49
; 
32'd34123: dataIn1 = 32'd50
; 
32'd34124: dataIn1 = 32'd51
; 
32'd34125: dataIn1 = 32'd52
; 
32'd34126: dataIn1 = 32'd53
; 
32'd34127: dataIn1 = 32'd55
; 
32'd34128: dataIn1 = 32'd56
; 
32'd34129: dataIn1 = 32'd58
; 
32'd34130: dataIn1 = 32'd59
; 
32'd34131: dataIn1 = 32'd60
; 
32'd34132: dataIn1 = 32'd62
; 
32'd34133: dataIn1 = 32'd0
; 
32'd34134: dataIn1 = 32'd1
; 
32'd34135: dataIn1 = 32'd2
; 
32'd34136: dataIn1 = 32'd3
; 
32'd34137: dataIn1 = 32'd6
; 
32'd34138: dataIn1 = 32'd7
; 
32'd34139: dataIn1 = 32'd8
; 
32'd34140: dataIn1 = 32'd9
; 
32'd34141: dataIn1 = 32'd14
; 
32'd34142: dataIn1 = 32'd17
; 
32'd34143: dataIn1 = 32'd18
; 
32'd34144: dataIn1 = 32'd23
; 
32'd34145: dataIn1 = 32'd24
; 
32'd34146: dataIn1 = 32'd25
; 
32'd34147: dataIn1 = 32'd26
; 
32'd34148: dataIn1 = 32'd27
; 
32'd34149: dataIn1 = 32'd31
; 
32'd34150: dataIn1 = 32'd32
; 
32'd34151: dataIn1 = 32'd34
; 
32'd34152: dataIn1 = 32'd35
; 
32'd34153: dataIn1 = 32'd36
; 
32'd34154: dataIn1 = 32'd38
; 
32'd34155: dataIn1 = 32'd39
; 
32'd34156: dataIn1 = 32'd40
; 
32'd34157: dataIn1 = 32'd41
; 
32'd34158: dataIn1 = 32'd42
; 
32'd34159: dataIn1 = 32'd43
; 
32'd34160: dataIn1 = 32'd44
; 
32'd34161: dataIn1 = 32'd46
; 
32'd34162: dataIn1 = 32'd47
; 
32'd34163: dataIn1 = 32'd48
; 
32'd34164: dataIn1 = 32'd49
; 
32'd34165: dataIn1 = 32'd50
; 
32'd34166: dataIn1 = 32'd51
; 
32'd34167: dataIn1 = 32'd52
; 
32'd34168: dataIn1 = 32'd53
; 
32'd34169: dataIn1 = 32'd55
; 
32'd34170: dataIn1 = 32'd56
; 
32'd34171: dataIn1 = 32'd57
; 
32'd34172: dataIn1 = 32'd58
; 
32'd34173: dataIn1 = 32'd61
; 
32'd34174: dataIn1 = 32'd62
; 
32'd34175: dataIn1 = 32'd1
; 
32'd34176: dataIn1 = 32'd2
; 
32'd34177: dataIn1 = 32'd3
; 
32'd34178: dataIn1 = 32'd5
; 
32'd34179: dataIn1 = 32'd6
; 
32'd34180: dataIn1 = 32'd8
; 
32'd34181: dataIn1 = 32'd9
; 
32'd34182: dataIn1 = 32'd10
; 
32'd34183: dataIn1 = 32'd11
; 
32'd34184: dataIn1 = 32'd12
; 
32'd34185: dataIn1 = 32'd14
; 
32'd34186: dataIn1 = 32'd15
; 
32'd34187: dataIn1 = 32'd16
; 
32'd34188: dataIn1 = 32'd17
; 
32'd34189: dataIn1 = 32'd18
; 
32'd34190: dataIn1 = 32'd20
; 
32'd34191: dataIn1 = 32'd21
; 
32'd34192: dataIn1 = 32'd23
; 
32'd34193: dataIn1 = 32'd25
; 
32'd34194: dataIn1 = 32'd26
; 
32'd34195: dataIn1 = 32'd27
; 
32'd34196: dataIn1 = 32'd29
; 
32'd34197: dataIn1 = 32'd30
; 
32'd34198: dataIn1 = 32'd31
; 
32'd34199: dataIn1 = 32'd32
; 
32'd34200: dataIn1 = 32'd35
; 
32'd34201: dataIn1 = 32'd41
; 
32'd34202: dataIn1 = 32'd42
; 
32'd34203: dataIn1 = 32'd43
; 
32'd34204: dataIn1 = 32'd46
; 
32'd34205: dataIn1 = 32'd47
; 
32'd34206: dataIn1 = 32'd49
; 
32'd34207: dataIn1 = 32'd50
; 
32'd34208: dataIn1 = 32'd51
; 
32'd34209: dataIn1 = 32'd53
; 
32'd34210: dataIn1 = 32'd55
; 
32'd34211: dataIn1 = 32'd56
; 
32'd34212: dataIn1 = 32'd58
; 
32'd34213: dataIn1 = 32'd59
; 
32'd34214: dataIn1 = 32'd60
; 
32'd34215: dataIn1 = 32'd62
; 
32'd34216: dataIn1 = 32'd63
; 
32'd34217: dataIn1 = 32'd1
; 
32'd34218: dataIn1 = 32'd4
; 
32'd34219: dataIn1 = 32'd5
; 
32'd34220: dataIn1 = 32'd6
; 
32'd34221: dataIn1 = 32'd8
; 
32'd34222: dataIn1 = 32'd11
; 
32'd34223: dataIn1 = 32'd12
; 
32'd34224: dataIn1 = 32'd14
; 
32'd34225: dataIn1 = 32'd15
; 
32'd34226: dataIn1 = 32'd16
; 
32'd34227: dataIn1 = 32'd18
; 
32'd34228: dataIn1 = 32'd21
; 
32'd34229: dataIn1 = 32'd22
; 
32'd34230: dataIn1 = 32'd23
; 
32'd34231: dataIn1 = 32'd24
; 
32'd34232: dataIn1 = 32'd25
; 
32'd34233: dataIn1 = 32'd26
; 
32'd34234: dataIn1 = 32'd28
; 
32'd34235: dataIn1 = 32'd29
; 
32'd34236: dataIn1 = 32'd31
; 
32'd34237: dataIn1 = 32'd32
; 
32'd34238: dataIn1 = 32'd34
; 
32'd34239: dataIn1 = 32'd35
; 
32'd34240: dataIn1 = 32'd36
; 
32'd34241: dataIn1 = 32'd39
; 
32'd34242: dataIn1 = 32'd40
; 
32'd34243: dataIn1 = 32'd41
; 
32'd34244: dataIn1 = 32'd42
; 
32'd34245: dataIn1 = 32'd43
; 
32'd34246: dataIn1 = 32'd44
; 
32'd34247: dataIn1 = 32'd45
; 
32'd34248: dataIn1 = 32'd47
; 
32'd34249: dataIn1 = 32'd50
; 
32'd34250: dataIn1 = 32'd52
; 
32'd34251: dataIn1 = 32'd53
; 
32'd34252: dataIn1 = 32'd55
; 
32'd34253: dataIn1 = 32'd56
; 
32'd34254: dataIn1 = 32'd57
; 
32'd34255: dataIn1 = 32'd60
; 
32'd34256: dataIn1 = 32'd61
; 
32'd34257: dataIn1 = 32'd0
; 
32'd34258: dataIn1 = 32'd1
; 
32'd34259: dataIn1 = 32'd2
; 
32'd34260: dataIn1 = 32'd3
; 
32'd34261: dataIn1 = 32'd6
; 
32'd34262: dataIn1 = 32'd7
; 
32'd34263: dataIn1 = 32'd8
; 
32'd34264: dataIn1 = 32'd9
; 
32'd34265: dataIn1 = 32'd11
; 
32'd34266: dataIn1 = 32'd12
; 
32'd34267: dataIn1 = 32'd14
; 
32'd34268: dataIn1 = 32'd15
; 
32'd34269: dataIn1 = 32'd16
; 
32'd34270: dataIn1 = 32'd17
; 
32'd34271: dataIn1 = 32'd19
; 
32'd34272: dataIn1 = 32'd20
; 
32'd34273: dataIn1 = 32'd23
; 
32'd34274: dataIn1 = 32'd25
; 
32'd34275: dataIn1 = 32'd27
; 
32'd34276: dataIn1 = 32'd28
; 
32'd34277: dataIn1 = 32'd30
; 
32'd34278: dataIn1 = 32'd31
; 
32'd34279: dataIn1 = 32'd33
; 
32'd34280: dataIn1 = 32'd34
; 
32'd34281: dataIn1 = 32'd36
; 
32'd34282: dataIn1 = 32'd38
; 
32'd34283: dataIn1 = 32'd39
; 
32'd34284: dataIn1 = 32'd40
; 
32'd34285: dataIn1 = 32'd43
; 
32'd34286: dataIn1 = 32'd45
; 
32'd34287: dataIn1 = 32'd46
; 
32'd34288: dataIn1 = 32'd47
; 
32'd34289: dataIn1 = 32'd48
; 
32'd34290: dataIn1 = 32'd49
; 
32'd34291: dataIn1 = 32'd50
; 
32'd34292: dataIn1 = 32'd52
; 
32'd34293: dataIn1 = 32'd53
; 
32'd34294: dataIn1 = 32'd55
; 
32'd34295: dataIn1 = 32'd56
; 
32'd34296: dataIn1 = 32'd59
; 
32'd34297: dataIn1 = 32'd61
; 
32'd34298: dataIn1 = 32'd62
; 
32'd34299: dataIn1 = 32'd0
; 
32'd34300: dataIn1 = 32'd1
; 
32'd34301: dataIn1 = 32'd3
; 
32'd34302: dataIn1 = 32'd4
; 
32'd34303: dataIn1 = 32'd6
; 
32'd34304: dataIn1 = 32'd7
; 
32'd34305: dataIn1 = 32'd11
; 
32'd34306: dataIn1 = 32'd12
; 
32'd34307: dataIn1 = 32'd13
; 
32'd34308: dataIn1 = 32'd14
; 
32'd34309: dataIn1 = 32'd15
; 
32'd34310: dataIn1 = 32'd16
; 
32'd34311: dataIn1 = 32'd17
; 
32'd34312: dataIn1 = 32'd20
; 
32'd34313: dataIn1 = 32'd21
; 
32'd34314: dataIn1 = 32'd22
; 
32'd34315: dataIn1 = 32'd24
; 
32'd34316: dataIn1 = 32'd26
; 
32'd34317: dataIn1 = 32'd27
; 
32'd34318: dataIn1 = 32'd29
; 
32'd34319: dataIn1 = 32'd30
; 
32'd34320: dataIn1 = 32'd31
; 
32'd34321: dataIn1 = 32'd35
; 
32'd34322: dataIn1 = 32'd36
; 
32'd34323: dataIn1 = 32'd37
; 
32'd34324: dataIn1 = 32'd38
; 
32'd34325: dataIn1 = 32'd40
; 
32'd34326: dataIn1 = 32'd42
; 
32'd34327: dataIn1 = 32'd44
; 
32'd34328: dataIn1 = 32'd45
; 
32'd34329: dataIn1 = 32'd46
; 
32'd34330: dataIn1 = 32'd47
; 
32'd34331: dataIn1 = 32'd48
; 
32'd34332: dataIn1 = 32'd51
; 
32'd34333: dataIn1 = 32'd53
; 
32'd34334: dataIn1 = 32'd55
; 
32'd34335: dataIn1 = 32'd56
; 
32'd34336: dataIn1 = 32'd57
; 
32'd34337: dataIn1 = 32'd58
; 
32'd34338: dataIn1 = 32'd59
; 
32'd34339: dataIn1 = 32'd62
; 
32'd34340: dataIn1 = 32'd63
; 
32'd34341: dataIn1 = 32'd0
; 
32'd34342: dataIn1 = 32'd1
; 
32'd34343: dataIn1 = 32'd2
; 
32'd34344: dataIn1 = 32'd4
; 
32'd34345: dataIn1 = 32'd5
; 
32'd34346: dataIn1 = 32'd6
; 
32'd34347: dataIn1 = 32'd8
; 
32'd34348: dataIn1 = 32'd9
; 
32'd34349: dataIn1 = 32'd10
; 
32'd34350: dataIn1 = 32'd13
; 
32'd34351: dataIn1 = 32'd14
; 
32'd34352: dataIn1 = 32'd15
; 
32'd34353: dataIn1 = 32'd21
; 
32'd34354: dataIn1 = 32'd23
; 
32'd34355: dataIn1 = 32'd24
; 
32'd34356: dataIn1 = 32'd25
; 
32'd34357: dataIn1 = 32'd28
; 
32'd34358: dataIn1 = 32'd29
; 
32'd34359: dataIn1 = 32'd30
; 
32'd34360: dataIn1 = 32'd32
; 
32'd34361: dataIn1 = 32'd33
; 
32'd34362: dataIn1 = 32'd34
; 
32'd34363: dataIn1 = 32'd37
; 
32'd34364: dataIn1 = 32'd38
; 
32'd34365: dataIn1 = 32'd39
; 
32'd34366: dataIn1 = 32'd40
; 
32'd34367: dataIn1 = 32'd41
; 
32'd34368: dataIn1 = 32'd43
; 
32'd34369: dataIn1 = 32'd44
; 
32'd34370: dataIn1 = 32'd47
; 
32'd34371: dataIn1 = 32'd48
; 
32'd34372: dataIn1 = 32'd49
; 
32'd34373: dataIn1 = 32'd51
; 
32'd34374: dataIn1 = 32'd52
; 
32'd34375: dataIn1 = 32'd53
; 
32'd34376: dataIn1 = 32'd54
; 
32'd34377: dataIn1 = 32'd56
; 
32'd34378: dataIn1 = 32'd57
; 
32'd34379: dataIn1 = 32'd58
; 
32'd34380: dataIn1 = 32'd59
; 
32'd34381: dataIn1 = 32'd60
; 
32'd34382: dataIn1 = 32'd61
; 
32'd34383: dataIn1 = 32'd62
; 
32'd34384: dataIn1 = 32'd63
; 
32'd34385: dataIn1 = 32'd0
; 
32'd34386: dataIn1 = 32'd1
; 
32'd34387: dataIn1 = 32'd2
; 
32'd34388: dataIn1 = 32'd3
; 
32'd34389: dataIn1 = 32'd4
; 
32'd34390: dataIn1 = 32'd7
; 
32'd34391: dataIn1 = 32'd11
; 
32'd34392: dataIn1 = 32'd12
; 
32'd34393: dataIn1 = 32'd13
; 
32'd34394: dataIn1 = 32'd14
; 
32'd34395: dataIn1 = 32'd15
; 
32'd34396: dataIn1 = 32'd16
; 
32'd34397: dataIn1 = 32'd17
; 
32'd34398: dataIn1 = 32'd19
; 
32'd34399: dataIn1 = 32'd20
; 
32'd34400: dataIn1 = 32'd21
; 
32'd34401: dataIn1 = 32'd22
; 
32'd34402: dataIn1 = 32'd23
; 
32'd34403: dataIn1 = 32'd24
; 
32'd34404: dataIn1 = 32'd25
; 
32'd34405: dataIn1 = 32'd27
; 
32'd34406: dataIn1 = 32'd28
; 
32'd34407: dataIn1 = 32'd30
; 
32'd34408: dataIn1 = 32'd31
; 
32'd34409: dataIn1 = 32'd32
; 
32'd34410: dataIn1 = 32'd33
; 
32'd34411: dataIn1 = 32'd37
; 
32'd34412: dataIn1 = 32'd38
; 
32'd34413: dataIn1 = 32'd42
; 
32'd34414: dataIn1 = 32'd44
; 
32'd34415: dataIn1 = 32'd46
; 
32'd34416: dataIn1 = 32'd47
; 
32'd34417: dataIn1 = 32'd48
; 
32'd34418: dataIn1 = 32'd49
; 
32'd34419: dataIn1 = 32'd50
; 
32'd34420: dataIn1 = 32'd51
; 
32'd34421: dataIn1 = 32'd52
; 
32'd34422: dataIn1 = 32'd54
; 
32'd34423: dataIn1 = 32'd55
; 
32'd34424: dataIn1 = 32'd56
; 
32'd34425: dataIn1 = 32'd57
; 
32'd34426: dataIn1 = 32'd62
; 
32'd34427: dataIn1 = 32'd63
; 
32'd34428: dataIn1 = 32'd0
; 
32'd34429: dataIn1 = 32'd1
; 
32'd34430: dataIn1 = 32'd3
; 
32'd34431: dataIn1 = 32'd4
; 
32'd34432: dataIn1 = 32'd6
; 
32'd34433: dataIn1 = 32'd7
; 
32'd34434: dataIn1 = 32'd8
; 
32'd34435: dataIn1 = 32'd9
; 
32'd34436: dataIn1 = 32'd10
; 
32'd34437: dataIn1 = 32'd12
; 
32'd34438: dataIn1 = 32'd16
; 
32'd34439: dataIn1 = 32'd18
; 
32'd34440: dataIn1 = 32'd23
; 
32'd34441: dataIn1 = 32'd24
; 
32'd34442: dataIn1 = 32'd25
; 
32'd34443: dataIn1 = 32'd26
; 
32'd34444: dataIn1 = 32'd27
; 
32'd34445: dataIn1 = 32'd28
; 
32'd34446: dataIn1 = 32'd33
; 
32'd34447: dataIn1 = 32'd34
; 
32'd34448: dataIn1 = 32'd35
; 
32'd34449: dataIn1 = 32'd36
; 
32'd34450: dataIn1 = 32'd37
; 
32'd34451: dataIn1 = 32'd38
; 
32'd34452: dataIn1 = 32'd40
; 
32'd34453: dataIn1 = 32'd41
; 
32'd34454: dataIn1 = 32'd42
; 
32'd34455: dataIn1 = 32'd44
; 
32'd34456: dataIn1 = 32'd45
; 
32'd34457: dataIn1 = 32'd46
; 
32'd34458: dataIn1 = 32'd47
; 
32'd34459: dataIn1 = 32'd49
; 
32'd34460: dataIn1 = 32'd50
; 
32'd34461: dataIn1 = 32'd51
; 
32'd34462: dataIn1 = 32'd52
; 
32'd34463: dataIn1 = 32'd53
; 
32'd34464: dataIn1 = 32'd54
; 
32'd34465: dataIn1 = 32'd55
; 
32'd34466: dataIn1 = 32'd58
; 
32'd34467: dataIn1 = 32'd60
; 
32'd34468: dataIn1 = 32'd63
; 
32'd34469: dataIn1 = 32'd0
; 
32'd34470: dataIn1 = 32'd1
; 
32'd34471: dataIn1 = 32'd2
; 
32'd34472: dataIn1 = 32'd4
; 
32'd34473: dataIn1 = 32'd5
; 
32'd34474: dataIn1 = 32'd6
; 
32'd34475: dataIn1 = 32'd8
; 
32'd34476: dataIn1 = 32'd9
; 
32'd34477: dataIn1 = 32'd10
; 
32'd34478: dataIn1 = 32'd11
; 
32'd34479: dataIn1 = 32'd12
; 
32'd34480: dataIn1 = 32'd13
; 
32'd34481: dataIn1 = 32'd14
; 
32'd34482: dataIn1 = 32'd15
; 
32'd34483: dataIn1 = 32'd16
; 
32'd34484: dataIn1 = 32'd17
; 
32'd34485: dataIn1 = 32'd18
; 
32'd34486: dataIn1 = 32'd19
; 
32'd34487: dataIn1 = 32'd20
; 
32'd34488: dataIn1 = 32'd21
; 
32'd34489: dataIn1 = 32'd22
; 
32'd34490: dataIn1 = 32'd23
; 
32'd34491: dataIn1 = 32'd24
; 
32'd34492: dataIn1 = 32'd25
; 
32'd34493: dataIn1 = 32'd26
; 
32'd34494: dataIn1 = 32'd27
; 
32'd34495: dataIn1 = 32'd28
; 
32'd34496: dataIn1 = 32'd29
; 
32'd34497: dataIn1 = 32'd30
; 
32'd34498: dataIn1 = 32'd31
; 
32'd34499: dataIn1 = 32'd32
; 
32'd34500: dataIn1 = 32'd36
; 
32'd34501: dataIn1 = 32'd37
; 
32'd34502: dataIn1 = 32'd38
; 
32'd34503: dataIn1 = 32'd39
; 
32'd34504: dataIn1 = 32'd40
; 
32'd34505: dataIn1 = 32'd42
; 
32'd34506: dataIn1 = 32'd43
; 
32'd34507: dataIn1 = 32'd44
; 
32'd34508: dataIn1 = 32'd46
; 
32'd34509: dataIn1 = 32'd47
; 
32'd34510: dataIn1 = 32'd49
; 
32'd34511: dataIn1 = 32'd50
; 
32'd34512: dataIn1 = 32'd51
; 
32'd34513: dataIn1 = 32'd52
; 
32'd34514: dataIn1 = 32'd53
; 
32'd34515: dataIn1 = 32'd54
; 
32'd34516: dataIn1 = 32'd55
; 
32'd34517: dataIn1 = 32'd57
; 
32'd34518: dataIn1 = 32'd62
; 
32'd34519: dataIn1 = 32'd63
; 
32'd34520: dataIn1 = 32'd0
; 
32'd34521: dataIn1 = 32'd3
; 
32'd34522: dataIn1 = 32'd4
; 
32'd34523: dataIn1 = 32'd5
; 
32'd34524: dataIn1 = 32'd6
; 
32'd34525: dataIn1 = 32'd7
; 
32'd34526: dataIn1 = 32'd9
; 
32'd34527: dataIn1 = 32'd10
; 
32'd34528: dataIn1 = 32'd11
; 
32'd34529: dataIn1 = 32'd18
; 
32'd34530: dataIn1 = 32'd19
; 
32'd34531: dataIn1 = 32'd20
; 
32'd34532: dataIn1 = 32'd21
; 
32'd34533: dataIn1 = 32'd22
; 
32'd34534: dataIn1 = 32'd23
; 
32'd34535: dataIn1 = 32'd28
; 
32'd34536: dataIn1 = 32'd29
; 
32'd34537: dataIn1 = 32'd30
; 
32'd34538: dataIn1 = 32'd31
; 
32'd34539: dataIn1 = 32'd34
; 
32'd34540: dataIn1 = 32'd35
; 
32'd34541: dataIn1 = 32'd38
; 
32'd34542: dataIn1 = 32'd39
; 
32'd34543: dataIn1 = 32'd40
; 
32'd34544: dataIn1 = 32'd43
; 
32'd34545: dataIn1 = 32'd46
; 
32'd34546: dataIn1 = 32'd47
; 
32'd34547: dataIn1 = 32'd48
; 
32'd34548: dataIn1 = 32'd51
; 
32'd34549: dataIn1 = 32'd52
; 
32'd34550: dataIn1 = 32'd53
; 
32'd34551: dataIn1 = 32'd54
; 
32'd34552: dataIn1 = 32'd57
; 
32'd34553: dataIn1 = 32'd58
; 
32'd34554: dataIn1 = 32'd59
; 
32'd34555: dataIn1 = 32'd61
; 
32'd34556: dataIn1 = 32'd63
; 
32'd34557: dataIn1 = 32'd1
; 
32'd34558: dataIn1 = 32'd2
; 
32'd34559: dataIn1 = 32'd3
; 
32'd34560: dataIn1 = 32'd4
; 
32'd34561: dataIn1 = 32'd5
; 
32'd34562: dataIn1 = 32'd6
; 
32'd34563: dataIn1 = 32'd8
; 
32'd34564: dataIn1 = 32'd9
; 
32'd34565: dataIn1 = 32'd10
; 
32'd34566: dataIn1 = 32'd11
; 
32'd34567: dataIn1 = 32'd12
; 
32'd34568: dataIn1 = 32'd14
; 
32'd34569: dataIn1 = 32'd15
; 
32'd34570: dataIn1 = 32'd17
; 
32'd34571: dataIn1 = 32'd18
; 
32'd34572: dataIn1 = 32'd19
; 
32'd34573: dataIn1 = 32'd20
; 
32'd34574: dataIn1 = 32'd22
; 
32'd34575: dataIn1 = 32'd24
; 
32'd34576: dataIn1 = 32'd26
; 
32'd34577: dataIn1 = 32'd27
; 
32'd34578: dataIn1 = 32'd29
; 
32'd34579: dataIn1 = 32'd34
; 
32'd34580: dataIn1 = 32'd35
; 
32'd34581: dataIn1 = 32'd36
; 
32'd34582: dataIn1 = 32'd38
; 
32'd34583: dataIn1 = 32'd39
; 
32'd34584: dataIn1 = 32'd41
; 
32'd34585: dataIn1 = 32'd44
; 
32'd34586: dataIn1 = 32'd45
; 
32'd34587: dataIn1 = 32'd47
; 
32'd34588: dataIn1 = 32'd50
; 
32'd34589: dataIn1 = 32'd52
; 
32'd34590: dataIn1 = 32'd53
; 
32'd34591: dataIn1 = 32'd54
; 
32'd34592: dataIn1 = 32'd56
; 
32'd34593: dataIn1 = 32'd57
; 
32'd34594: dataIn1 = 32'd58
; 
32'd34595: dataIn1 = 32'd59
; 
32'd34596: dataIn1 = 32'd62
; 
32'd34597: dataIn1 = 32'd0
; 
32'd34598: dataIn1 = 32'd1
; 
32'd34599: dataIn1 = 32'd2
; 
32'd34600: dataIn1 = 32'd5
; 
32'd34601: dataIn1 = 32'd7
; 
32'd34602: dataIn1 = 32'd9
; 
32'd34603: dataIn1 = 32'd10
; 
32'd34604: dataIn1 = 32'd11
; 
32'd34605: dataIn1 = 32'd12
; 
32'd34606: dataIn1 = 32'd13
; 
32'd34607: dataIn1 = 32'd14
; 
32'd34608: dataIn1 = 32'd15
; 
32'd34609: dataIn1 = 32'd16
; 
32'd34610: dataIn1 = 32'd17
; 
32'd34611: dataIn1 = 32'd18
; 
32'd34612: dataIn1 = 32'd21
; 
32'd34613: dataIn1 = 32'd22
; 
32'd34614: dataIn1 = 32'd24
; 
32'd34615: dataIn1 = 32'd25
; 
32'd34616: dataIn1 = 32'd26
; 
32'd34617: dataIn1 = 32'd27
; 
32'd34618: dataIn1 = 32'd28
; 
32'd34619: dataIn1 = 32'd29
; 
32'd34620: dataIn1 = 32'd30
; 
32'd34621: dataIn1 = 32'd31
; 
32'd34622: dataIn1 = 32'd32
; 
32'd34623: dataIn1 = 32'd33
; 
32'd34624: dataIn1 = 32'd35
; 
32'd34625: dataIn1 = 32'd36
; 
32'd34626: dataIn1 = 32'd37
; 
32'd34627: dataIn1 = 32'd40
; 
32'd34628: dataIn1 = 32'd41
; 
32'd34629: dataIn1 = 32'd42
; 
32'd34630: dataIn1 = 32'd43
; 
32'd34631: dataIn1 = 32'd45
; 
32'd34632: dataIn1 = 32'd48
; 
32'd34633: dataIn1 = 32'd49
; 
32'd34634: dataIn1 = 32'd50
; 
32'd34635: dataIn1 = 32'd51
; 
32'd34636: dataIn1 = 32'd52
; 
32'd34637: dataIn1 = 32'd54
; 
32'd34638: dataIn1 = 32'd55
; 
32'd34639: dataIn1 = 32'd56
; 
32'd34640: dataIn1 = 32'd58
; 
32'd34641: dataIn1 = 32'd60
; 
32'd34642: dataIn1 = 32'd61
; 
32'd34643: dataIn1 = 32'd63
; 
32'd34644: dataIn1 = 32'd1
; 
32'd34645: dataIn1 = 32'd2
; 
32'd34646: dataIn1 = 32'd3
; 
32'd34647: dataIn1 = 32'd4
; 
32'd34648: dataIn1 = 32'd5
; 
32'd34649: dataIn1 = 32'd6
; 
32'd34650: dataIn1 = 32'd7
; 
32'd34651: dataIn1 = 32'd8
; 
32'd34652: dataIn1 = 32'd9
; 
32'd34653: dataIn1 = 32'd12
; 
32'd34654: dataIn1 = 32'd15
; 
32'd34655: dataIn1 = 32'd21
; 
32'd34656: dataIn1 = 32'd23
; 
32'd34657: dataIn1 = 32'd24
; 
32'd34658: dataIn1 = 32'd26
; 
32'd34659: dataIn1 = 32'd27
; 
32'd34660: dataIn1 = 32'd28
; 
32'd34661: dataIn1 = 32'd30
; 
32'd34662: dataIn1 = 32'd34
; 
32'd34663: dataIn1 = 32'd35
; 
32'd34664: dataIn1 = 32'd36
; 
32'd34665: dataIn1 = 32'd37
; 
32'd34666: dataIn1 = 32'd39
; 
32'd34667: dataIn1 = 32'd42
; 
32'd34668: dataIn1 = 32'd44
; 
32'd34669: dataIn1 = 32'd45
; 
32'd34670: dataIn1 = 32'd46
; 
32'd34671: dataIn1 = 32'd47
; 
32'd34672: dataIn1 = 32'd49
; 
32'd34673: dataIn1 = 32'd50
; 
32'd34674: dataIn1 = 32'd51
; 
32'd34675: dataIn1 = 32'd52
; 
32'd34676: dataIn1 = 32'd53
; 
32'd34677: dataIn1 = 32'd54
; 
32'd34678: dataIn1 = 32'd55
; 
32'd34679: dataIn1 = 32'd56
; 
32'd34680: dataIn1 = 32'd58
; 
32'd34681: dataIn1 = 32'd59
; 
32'd34682: dataIn1 = 32'd61
; 
32'd34683: dataIn1 = 32'd62
; 
32'd34684: dataIn1 = 32'd63
; 
32'd34685: dataIn1 = 32'd0
; 
32'd34686: dataIn1 = 32'd1
; 
32'd34687: dataIn1 = 32'd2
; 
32'd34688: dataIn1 = 32'd4
; 
32'd34689: dataIn1 = 32'd7
; 
32'd34690: dataIn1 = 32'd9
; 
32'd34691: dataIn1 = 32'd11
; 
32'd34692: dataIn1 = 32'd13
; 
32'd34693: dataIn1 = 32'd15
; 
32'd34694: dataIn1 = 32'd17
; 
32'd34695: dataIn1 = 32'd18
; 
32'd34696: dataIn1 = 32'd19
; 
32'd34697: dataIn1 = 32'd21
; 
32'd34698: dataIn1 = 32'd22
; 
32'd34699: dataIn1 = 32'd23
; 
32'd34700: dataIn1 = 32'd24
; 
32'd34701: dataIn1 = 32'd25
; 
32'd34702: dataIn1 = 32'd27
; 
32'd34703: dataIn1 = 32'd29
; 
32'd34704: dataIn1 = 32'd30
; 
32'd34705: dataIn1 = 32'd32
; 
32'd34706: dataIn1 = 32'd33
; 
32'd34707: dataIn1 = 32'd34
; 
32'd34708: dataIn1 = 32'd35
; 
32'd34709: dataIn1 = 32'd37
; 
32'd34710: dataIn1 = 32'd38
; 
32'd34711: dataIn1 = 32'd39
; 
32'd34712: dataIn1 = 32'd41
; 
32'd34713: dataIn1 = 32'd42
; 
32'd34714: dataIn1 = 32'd43
; 
32'd34715: dataIn1 = 32'd45
; 
32'd34716: dataIn1 = 32'd50
; 
32'd34717: dataIn1 = 32'd51
; 
32'd34718: dataIn1 = 32'd53
; 
32'd34719: dataIn1 = 32'd55
; 
32'd34720: dataIn1 = 32'd56
; 
32'd34721: dataIn1 = 32'd57
; 
32'd34722: dataIn1 = 32'd58
; 
32'd34723: dataIn1 = 32'd59
; 
32'd34724: dataIn1 = 32'd60
; 
32'd34725: dataIn1 = 32'd62
; 
32'd34726: dataIn1 = 32'd63
; 
32'd34727: dataIn1 = 32'd1
; 
32'd34728: dataIn1 = 32'd5
; 
32'd34729: dataIn1 = 32'd6
; 
32'd34730: dataIn1 = 32'd7
; 
32'd34731: dataIn1 = 32'd8
; 
32'd34732: dataIn1 = 32'd9
; 
32'd34733: dataIn1 = 32'd11
; 
32'd34734: dataIn1 = 32'd12
; 
32'd34735: dataIn1 = 32'd13
; 
32'd34736: dataIn1 = 32'd14
; 
32'd34737: dataIn1 = 32'd16
; 
32'd34738: dataIn1 = 32'd17
; 
32'd34739: dataIn1 = 32'd19
; 
32'd34740: dataIn1 = 32'd20
; 
32'd34741: dataIn1 = 32'd21
; 
32'd34742: dataIn1 = 32'd22
; 
32'd34743: dataIn1 = 32'd24
; 
32'd34744: dataIn1 = 32'd26
; 
32'd34745: dataIn1 = 32'd28
; 
32'd34746: dataIn1 = 32'd30
; 
32'd34747: dataIn1 = 32'd31
; 
32'd34748: dataIn1 = 32'd32
; 
32'd34749: dataIn1 = 32'd33
; 
32'd34750: dataIn1 = 32'd35
; 
32'd34751: dataIn1 = 32'd38
; 
32'd34752: dataIn1 = 32'd39
; 
32'd34753: dataIn1 = 32'd40
; 
32'd34754: dataIn1 = 32'd41
; 
32'd34755: dataIn1 = 32'd42
; 
32'd34756: dataIn1 = 32'd43
; 
32'd34757: dataIn1 = 32'd44
; 
32'd34758: dataIn1 = 32'd45
; 
32'd34759: dataIn1 = 32'd46
; 
32'd34760: dataIn1 = 32'd47
; 
32'd34761: dataIn1 = 32'd48
; 
32'd34762: dataIn1 = 32'd50
; 
32'd34763: dataIn1 = 32'd52
; 
32'd34764: dataIn1 = 32'd54
; 
32'd34765: dataIn1 = 32'd56
; 
32'd34766: dataIn1 = 32'd57
; 
32'd34767: dataIn1 = 32'd59
; 
32'd34768: dataIn1 = 32'd60
; 
32'd34769: dataIn1 = 32'd62
; 
32'd34770: dataIn1 = 32'd63
; 
32'd34771: dataIn1 = 32'd0
; 
32'd34772: dataIn1 = 32'd2
; 
32'd34773: dataIn1 = 32'd3
; 
32'd34774: dataIn1 = 32'd4
; 
32'd34775: dataIn1 = 32'd5
; 
32'd34776: dataIn1 = 32'd9
; 
32'd34777: dataIn1 = 32'd10
; 
32'd34778: dataIn1 = 32'd12
; 
32'd34779: dataIn1 = 32'd14
; 
32'd34780: dataIn1 = 32'd16
; 
32'd34781: dataIn1 = 32'd19
; 
32'd34782: dataIn1 = 32'd20
; 
32'd34783: dataIn1 = 32'd21
; 
32'd34784: dataIn1 = 32'd23
; 
32'd34785: dataIn1 = 32'd24
; 
32'd34786: dataIn1 = 32'd28
; 
32'd34787: dataIn1 = 32'd30
; 
32'd34788: dataIn1 = 32'd32
; 
32'd34789: dataIn1 = 32'd33
; 
32'd34790: dataIn1 = 32'd34
; 
32'd34791: dataIn1 = 32'd36
; 
32'd34792: dataIn1 = 32'd37
; 
32'd34793: dataIn1 = 32'd38
; 
32'd34794: dataIn1 = 32'd40
; 
32'd34795: dataIn1 = 32'd42
; 
32'd34796: dataIn1 = 32'd46
; 
32'd34797: dataIn1 = 32'd48
; 
32'd34798: dataIn1 = 32'd49
; 
32'd34799: dataIn1 = 32'd51
; 
32'd34800: dataIn1 = 32'd53
; 
32'd34801: dataIn1 = 32'd54
; 
32'd34802: dataIn1 = 32'd55
; 
32'd34803: dataIn1 = 32'd56
; 
32'd34804: dataIn1 = 32'd57
; 
32'd34805: dataIn1 = 32'd59
; 
32'd34806: dataIn1 = 32'd62
; 
32'd34807: dataIn1 = 32'd63
; 
32'd34808: dataIn1 = 32'd; 
32'd34809: dataIn1 = 32'd; 
32'd34810: dataIn1 = 32'd; 
32'd34811: dataIn1 = 32'd; 
32'd34812: dataIn1 = 32'd; 
32'd34813: dataIn1 = 32'd; 
32'd34814: dataIn1 = 32'd; 
32'd34815: dataIn1 = 32'd; 
32'd34816: dataIn1 = 32'd; 
32'd34817: dataIn1 = 32'd; 
32'd34818: dataIn1 = 32'd; 
32'd34819: dataIn1 = 32'd; 
32'd34820: dataIn1 = 32'd; 
32'd34821: dataIn1 = 32'd; 
32'd34822: dataIn1 = 32'd; 
32'd34823: dataIn1 = 32'd; 
32'd34824: dataIn1 = 32'd; 
32'd34825: dataIn1 = 32'd; 
32'd34826: dataIn1 = 32'd; 
32'd34827: dataIn1 = 32'd; 
32'd34828: dataIn1 = 32'd; 
32'd34829: dataIn1 = 32'd; 
32'd34830: dataIn1 = 32'd; 
32'd34831: dataIn1 = 32'd; 
32'd34832: dataIn1 = 32'd; 
32'd34833: dataIn1 = 32'd; 
32'd34834: dataIn1 = 32'd; 
32'd34835: dataIn1 = 32'd; 
32'd34836: dataIn1 = 32'd; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd4; 
32'd3: dataIn2 = 32'd20; 
32'd4: dataIn2 = 32'd90; 
32'd5: dataIn2 = 32'd0; 
32'd6: dataIn2 = 32'd22; 
32'd7: dataIn2 = 32'd2; 
32'd8: dataIn2 = 32'd81; 
32'd9: dataIn2 = 32'd1; 
32'd10: dataIn2 = 32'd77; 
32'd11: dataIn2 = 32'd70; 
32'd12: dataIn2 = 32'd24; 
32'd13: dataIn2 = 32'd41; 
32'd14: dataIn2 = 32'd60; 
32'd15: dataIn2 = 32'd20; 
32'd16: dataIn2 = 32'd44; 
32'd17: dataIn2 = 32'd55; 
32'd18: dataIn2 = 32'd31; 
32'd19: dataIn2 = 32'd71; 
32'd20: dataIn2 = 32'd21; 
32'd21: dataIn2 = 32'd38; 
32'd22: dataIn2 = 32'd15; 
32'd23: dataIn2 = 32'd2; 
32'd24: dataIn2 = 32'd51; 
32'd25: dataIn2 = 32'd56; 
32'd26: dataIn2 = 32'd94; 
32'd27: dataIn2 = 32'd64; 
32'd28: dataIn2 = 32'd53; 
32'd29: dataIn2 = 32'd16; 
32'd30: dataIn2 = 32'd75; 
32'd31: dataIn2 = 32'd61; 
32'd32: dataIn2 = 32'd88; 
32'd33: dataIn2 = 32'd0; 
32'd34: dataIn2 = 32'd2; 
32'd35: dataIn2 = 32'd88; 
32'd36: dataIn2 = 32'd60; 
32'd37: dataIn2 = 32'd93; 
32'd38: dataIn2 = 32'd51; 
32'd39: dataIn2 = 32'd55; 
32'd40: dataIn2 = 32'd78; 
32'd41: dataIn2 = 32'd27; 
32'd42: dataIn2 = 32'd67; 
32'd43: dataIn2 = 32'd47; 
32'd44: dataIn2 = 32'd66; 
32'd45: dataIn2 = 32'd12; 
32'd46: dataIn2 = 32'd63; 
32'd47: dataIn2 = 32'd94; 
32'd48: dataIn2 = 32'd1; 
32'd49: dataIn2 = 32'd23; 
32'd50: dataIn2 = 32'd99; 
32'd51: dataIn2 = 32'd18; 
32'd52: dataIn2 = 32'd35; 
32'd53: dataIn2 = 32'd1; 
32'd54: dataIn2 = 32'd11; 
32'd55: dataIn2 = 32'd71; 
32'd56: dataIn2 = 32'd93; 
32'd57: dataIn2 = 32'd62; 
32'd58: dataIn2 = 32'd41; 
32'd59: dataIn2 = 32'd72; 
32'd60: dataIn2 = 32'd94; 
32'd61: dataIn2 = 32'd87; 
32'd62: dataIn2 = 32'd20; 
32'd63: dataIn2 = 32'd88; 
32'd64: dataIn2 = 32'd3; 
32'd65: dataIn2 = 32'd25; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd330: dataIn2 = 32'd2; 
32'd331: dataIn2 = 32'd37; 
32'd332: dataIn2 = 32'd7; 
32'd333: dataIn2 = 32'd62; 
32'd334: dataIn2 = 32'd84; 
32'd335: dataIn2 = 32'd27; 
32'd336: dataIn2 = 32'd72; 
32'd337: dataIn2 = 32'd27; 
32'd338: dataIn2 = 32'd35; 
32'd339: dataIn2 = 32'd94; 
32'd340: dataIn2 = 32'd95; 
32'd341: dataIn2 = 32'd52; 
32'd342: dataIn2 = 32'd59; 
32'd343: dataIn2 = 32'd47; 
32'd344: dataIn2 = 32'd40; 
32'd345: dataIn2 = 32'd10; 
32'd346: dataIn2 = 32'd28; 
32'd347: dataIn2 = 32'd95; 
32'd348: dataIn2 = 32'd21; 
32'd349: dataIn2 = 32'd45; 
32'd350: dataIn2 = 32'd74; 
32'd351: dataIn2 = 32'd4; 
32'd352: dataIn2 = 32'd3; 
32'd353: dataIn2 = 32'd48; 
32'd354: dataIn2 = 32'd89; 
32'd355: dataIn2 = 32'd99; 
32'd356: dataIn2 = 32'd24; 
32'd357: dataIn2 = 32'd38; 
32'd358: dataIn2 = 32'd64; 
32'd359: dataIn2 = 32'd95; 
32'd360: dataIn2 = 32'd5; 
32'd361: dataIn2 = 32'd70; 
32'd362: dataIn2 = 32'd97; 
32'd363: dataIn2 = 32'd82; 
32'd364: dataIn2 = 32'd16; 
32'd365: dataIn2 = 32'd45; 
32'd366: dataIn2 = 32'd49; 
32'd367: dataIn2 = 32'd61; 
32'd368: dataIn2 = 32'd16; 
32'd369: dataIn2 = 32'd0; 
32'd370: dataIn2 = 32'd56; 
32'd371: dataIn2 = 32'd75; 
32'd372: dataIn2 = 32'd98; 
32'd373: dataIn2 = 32'd85; 
32'd374: dataIn2 = 32'd7; 
32'd375: dataIn2 = 32'd66; 
32'd376: dataIn2 = 32'd46; 
32'd377: dataIn2 = 32'd62; 
32'd378: dataIn2 = 32'd80; 
32'd379: dataIn2 = 32'd100; 
32'd380: dataIn2 = 32'd77; 
32'd381: dataIn2 = 32'd39; 
32'd382: dataIn2 = 32'd26; 
32'd383: dataIn2 = 32'd95; 
32'd384: dataIn2 = 32'd77; 
32'd385: dataIn2 = 32'd41; 
32'd386: dataIn2 = 32'd19; 
32'd387: dataIn2 = 32'd5; 
32'd388: dataIn2 = 32'd46; 
32'd389: dataIn2 = 32'd36; 
32'd390: dataIn2 = 32'd39; 
32'd391: dataIn2 = 32'd64; 
32'd392: dataIn2 = 32'd86; 
32'd393: dataIn2 = 32'd28; 
32'd394: dataIn2 = 32'd76; 
32'd395: dataIn2 = 32'd99; 
32'd396: dataIn2 = 32'd87; 
32'd397: dataIn2 = 32'd69; 
32'd398: dataIn2 = 32'd17; 
32'd399: dataIn2 = 32'd68; 
32'd400: dataIn2 = 32'd86; 
32'd401: dataIn2 = 32'd90; 
32'd402: dataIn2 = 32'd31; 
32'd403: dataIn2 = 32'd43; 
32'd404: dataIn2 = 32'd62; 
32'd405: dataIn2 = 32'd41; 
32'd406: dataIn2 = 32'd35; 
32'd407: dataIn2 = 32'd2; 
32'd408: dataIn2 = 32'd86; 
32'd409: dataIn2 = 32'd23; 
32'd410: dataIn2 = 32'd16; 
32'd411: dataIn2 = 32'd69; 
32'd412: dataIn2 = 32'd37; 
32'd413: dataIn2 = 32'd0; 
32'd414: dataIn2 = 32'd52; 
32'd415: dataIn2 = 32'd37; 
32'd416: dataIn2 = 32'd53; 
32'd417: dataIn2 = 32'd28; 
32'd418: dataIn2 = 32'd69; 
32'd419: dataIn2 = 32'd53; 
32'd420: dataIn2 = 32'd38; 
32'd421: dataIn2 = 32'd61; 
32'd422: dataIn2 = 32'd40; 
32'd423: dataIn2 = 32'd100; 
32'd424: dataIn2 = 32'd42; 
32'd425: dataIn2 = 32'd38; 
32'd426: dataIn2 = 32'd46; 
32'd427: dataIn2 = 32'd56; 
32'd428: dataIn2 = 32'd66; 
32'd429: dataIn2 = 32'd74; 
32'd430: dataIn2 = 32'd7; 
32'd431: dataIn2 = 32'd83; 
32'd432: dataIn2 = 32'd69; 
32'd433: dataIn2 = 32'd42; 
32'd434: dataIn2 = 32'd43; 
32'd435: dataIn2 = 32'd73; 
32'd436: dataIn2 = 32'd62; 
32'd437: dataIn2 = 32'd23; 
32'd438: dataIn2 = 32'd98; 
32'd439: dataIn2 = 32'd31; 
32'd440: dataIn2 = 32'd22; 
32'd441: dataIn2 = 32'd41; 
32'd442: dataIn2 = 32'd80; 
32'd443: dataIn2 = 32'd19; 
32'd444: dataIn2 = 32'd96; 
32'd445: dataIn2 = 32'd72; 
32'd446: dataIn2 = 32'd16; 
32'd447: dataIn2 = 32'd57; 
32'd448: dataIn2 = 32'd31; 
32'd449: dataIn2 = 32'd27; 
32'd450: dataIn2 = 32'd67; 
32'd451: dataIn2 = 32'd18; 
32'd452: dataIn2 = 32'd82; 
32'd453: dataIn2 = 32'd64; 
32'd454: dataIn2 = 32'd86; 
32'd455: dataIn2 = 32'd18; 
32'd456: dataIn2 = 32'd21; 
32'd457: dataIn2 = 32'd69; 
32'd458: dataIn2 = 32'd58; 
32'd459: dataIn2 = 32'd41; 
32'd460: dataIn2 = 32'd56; 
32'd461: dataIn2 = 32'd23; 
32'd462: dataIn2 = 32'd43; 
32'd463: dataIn2 = 32'd88; 
32'd464: dataIn2 = 32'd81; 
32'd465: dataIn2 = 32'd84; 
32'd466: dataIn2 = 32'd74; 
32'd467: dataIn2 = 32'd94; 
32'd468: dataIn2 = 32'd54; 
32'd469: dataIn2 = 32'd79; 
32'd470: dataIn2 = 32'd40; 
32'd471: dataIn2 = 32'd80; 
32'd472: dataIn2 = 32'd91; 
32'd473: dataIn2 = 32'd66; 
32'd474: dataIn2 = 32'd7; 
32'd475: dataIn2 = 32'd64; 
32'd476: dataIn2 = 32'd34; 
32'd477: dataIn2 = 32'd36; 
32'd478: dataIn2 = 32'd7; 
32'd479: dataIn2 = 32'd3; 
32'd480: dataIn2 = 32'd97; 
32'd481: dataIn2 = 32'd27; 
32'd482: dataIn2 = 32'd13; 
32'd483: dataIn2 = 32'd39; 
32'd484: dataIn2 = 32'd10; 
32'd485: dataIn2 = 32'd65; 
32'd486: dataIn2 = 32'd20; 
32'd487: dataIn2 = 32'd91; 
32'd488: dataIn2 = 32'd86; 
32'd489: dataIn2 = 32'd50; 
32'd490: dataIn2 = 32'd64; 
32'd491: dataIn2 = 32'd11; 
32'd492: dataIn2 = 32'd30; 
32'd493: dataIn2 = 32'd0; 
32'd494: dataIn2 = 32'd19; 
32'd495: dataIn2 = 32'd1; 
32'd496: dataIn2 = 32'd91; 
32'd497: dataIn2 = 32'd11; 
32'd498: dataIn2 = 32'd77; 
32'd499: dataIn2 = 32'd47; 
32'd500: dataIn2 = 32'd86; 
32'd501: dataIn2 = 32'd22; 
32'd502: dataIn2 = 32'd75; 
32'd503: dataIn2 = 32'd72; 
32'd504: dataIn2 = 32'd26; 
32'd505: dataIn2 = 32'd25; 
32'd506: dataIn2 = 32'd24; 
32'd507: dataIn2 = 32'd46; 
32'd508: dataIn2 = 32'd79; 
32'd509: dataIn2 = 32'd80; 
32'd510: dataIn2 = 32'd50; 
32'd511: dataIn2 = 32'd32; 
32'd512: dataIn2 = 32'd16; 
32'd513: dataIn2 = 32'd55; 
32'd514: dataIn2 = 32'd33; 
32'd515: dataIn2 = 32'd10; 
32'd516: dataIn2 = 32'd13; 
32'd517: dataIn2 = 32'd63; 
32'd518: dataIn2 = 32'd48; 
32'd519: dataIn2 = 32'd84; 
32'd520: dataIn2 = 32'd10; 
32'd521: dataIn2 = 32'd52; 
32'd522: dataIn2 = 32'd11; 
32'd523: dataIn2 = 32'd14; 
32'd524: dataIn2 = 32'd84; 
32'd525: dataIn2 = 32'd7; 
32'd526: dataIn2 = 32'd15; 
32'd527: dataIn2 = 32'd41; 
32'd528: dataIn2 = 32'd22; 
32'd529: dataIn2 = 32'd37; 
32'd530: dataIn2 = 32'd40; 
32'd531: dataIn2 = 32'd97; 
32'd532: dataIn2 = 32'd36; 
32'd533: dataIn2 = 32'd61; 
32'd534: dataIn2 = 32'd81; 
32'd535: dataIn2 = 32'd14; 
32'd536: dataIn2 = 32'd98; 
32'd537: dataIn2 = 32'd88; 
32'd538: dataIn2 = 32'd32; 
32'd539: dataIn2 = 32'd57; 
32'd540: dataIn2 = 32'd97; 
32'd541: dataIn2 = 32'd75; 
32'd542: dataIn2 = 32'd63; 
32'd543: dataIn2 = 32'd98; 
32'd544: dataIn2 = 32'd65; 
32'd545: dataIn2 = 32'd23; 
32'd546: dataIn2 = 32'd26; 
32'd547: dataIn2 = 32'd44; 
32'd548: dataIn2 = 32'd9; 
32'd549: dataIn2 = 32'd92; 
32'd550: dataIn2 = 32'd12; 
32'd551: dataIn2 = 32'd70; 
32'd552: dataIn2 = 32'd17; 
32'd553: dataIn2 = 32'd54; 
32'd554: dataIn2 = 32'd49; 
32'd555: dataIn2 = 32'd18; 
32'd556: dataIn2 = 32'd87; 
32'd557: dataIn2 = 32'd60; 
32'd558: dataIn2 = 32'd84; 
32'd559: dataIn2 = 32'd27; 
32'd560: dataIn2 = 32'd43; 
32'd561: dataIn2 = 32'd65; 
32'd562: dataIn2 = 32'd39; 
32'd563: dataIn2 = 32'd18; 
32'd564: dataIn2 = 32'd22; 
32'd565: dataIn2 = 32'd41; 
32'd566: dataIn2 = 32'd80; 
32'd567: dataIn2 = 32'd50; 
32'd568: dataIn2 = 32'd71; 
32'd569: dataIn2 = 32'd0; 
32'd570: dataIn2 = 32'd76; 
32'd571: dataIn2 = 32'd90; 
32'd572: dataIn2 = 32'd46; 
32'd573: dataIn2 = 32'd14; 
32'd574: dataIn2 = 32'd28; 
32'd575: dataIn2 = 32'd67; 
32'd576: dataIn2 = 32'd18; 
32'd577: dataIn2 = 32'd93; 
32'd578: dataIn2 = 32'd90; 
32'd579: dataIn2 = 32'd100; 
32'd580: dataIn2 = 32'd50; 
32'd581: dataIn2 = 32'd29; 
32'd582: dataIn2 = 32'd1; 
32'd583: dataIn2 = 32'd95; 
32'd584: dataIn2 = 32'd9; 
32'd585: dataIn2 = 32'd63; 
32'd586: dataIn2 = 32'd73; 
32'd587: dataIn2 = 32'd75; 
32'd588: dataIn2 = 32'd37; 
32'd589: dataIn2 = 32'd30; 
32'd590: dataIn2 = 32'd94; 
32'd591: dataIn2 = 32'd43; 
32'd592: dataIn2 = 32'd34; 
32'd593: dataIn2 = 32'd43; 
32'd594: dataIn2 = 32'd39; 
32'd595: dataIn2 = 32'd74; 
32'd596: dataIn2 = 32'd29; 
32'd597: dataIn2 = 32'd90; 
32'd598: dataIn2 = 32'd47; 
32'd599: dataIn2 = 32'd21; 
32'd600: dataIn2 = 32'd51; 
32'd601: dataIn2 = 32'd56; 
32'd602: dataIn2 = 32'd25; 
32'd603: dataIn2 = 32'd39; 
32'd604: dataIn2 = 32'd41; 
32'd605: dataIn2 = 32'd78; 
32'd606: dataIn2 = 32'd47; 
32'd607: dataIn2 = 32'd10; 
32'd608: dataIn2 = 32'd79; 
32'd609: dataIn2 = 32'd51; 
32'd610: dataIn2 = 32'd90; 
32'd611: dataIn2 = 32'd92; 
32'd612: dataIn2 = 32'd52; 
32'd613: dataIn2 = 32'd78; 
32'd614: dataIn2 = 32'd27; 
32'd615: dataIn2 = 32'd46; 
32'd616: dataIn2 = 32'd18; 
32'd617: dataIn2 = 32'd17; 
32'd618: dataIn2 = 32'd56; 
32'd619: dataIn2 = 32'd28; 
32'd620: dataIn2 = 32'd70; 
32'd621: dataIn2 = 32'd68; 
32'd622: dataIn2 = 32'd72; 
32'd623: dataIn2 = 32'd41; 
32'd624: dataIn2 = 32'd52; 
32'd625: dataIn2 = 32'd4; 
32'd626: dataIn2 = 32'd27; 
32'd627: dataIn2 = 32'd4; 
32'd628: dataIn2 = 32'd26; 
32'd629: dataIn2 = 32'd61; 
32'd630: dataIn2 = 32'd84; 
32'd631: dataIn2 = 32'd0; 
32'd632: dataIn2 = 32'd7; 
32'd633: dataIn2 = 32'd12; 
32'd634: dataIn2 = 32'd28; 
32'd635: dataIn2 = 32'd61; 
32'd636: dataIn2 = 32'd5; 
32'd637: dataIn2 = 32'd56; 
32'd638: dataIn2 = 32'd94; 
32'd639: dataIn2 = 32'd63; 
32'd640: dataIn2 = 32'd62; 
32'd641: dataIn2 = 32'd52; 
32'd642: dataIn2 = 32'd52; 
32'd643: dataIn2 = 32'd8; 
32'd644: dataIn2 = 32'd56; 
32'd645: dataIn2 = 32'd50; 
32'd646: dataIn2 = 32'd78; 
32'd647: dataIn2 = 32'd100; 
32'd648: dataIn2 = 32'd62; 
32'd649: dataIn2 = 32'd41; 
32'd650: dataIn2 = 32'd84; 
32'd651: dataIn2 = 32'd70; 
32'd652: dataIn2 = 32'd95; 
32'd653: dataIn2 = 32'd89; 
32'd654: dataIn2 = 32'd68; 
32'd655: dataIn2 = 32'd9; 
32'd656: dataIn2 = 32'd23; 
32'd657: dataIn2 = 32'd18; 
32'd658: dataIn2 = 32'd42; 
32'd659: dataIn2 = 32'd61; 
32'd660: dataIn2 = 32'd68; 
32'd661: dataIn2 = 32'd32; 
32'd662: dataIn2 = 32'd14; 
32'd663: dataIn2 = 32'd58; 
32'd664: dataIn2 = 32'd56; 
32'd665: dataIn2 = 32'd85; 
32'd666: dataIn2 = 32'd82; 
32'd667: dataIn2 = 32'd61; 
32'd668: dataIn2 = 32'd88; 
32'd669: dataIn2 = 32'd60; 
32'd670: dataIn2 = 32'd8; 
32'd671: dataIn2 = 32'd66; 
32'd672: dataIn2 = 32'd11; 
32'd673: dataIn2 = 32'd74; 
32'd674: dataIn2 = 32'd100; 
32'd675: dataIn2 = 32'd67; 
32'd676: dataIn2 = 32'd94; 
32'd677: dataIn2 = 32'd47; 
32'd678: dataIn2 = 32'd48; 
32'd679: dataIn2 = 32'd22; 
32'd680: dataIn2 = 32'd45; 
32'd681: dataIn2 = 32'd89; 
32'd682: dataIn2 = 32'd97; 
32'd683: dataIn2 = 32'd99; 
32'd684: dataIn2 = 32'd31; 
32'd685: dataIn2 = 32'd20; 
32'd686: dataIn2 = 32'd100; 
32'd687: dataIn2 = 32'd68; 
32'd688: dataIn2 = 32'd66; 
32'd689: dataIn2 = 32'd80; 
32'd690: dataIn2 = 32'd23; 
32'd691: dataIn2 = 32'd97; 
32'd692: dataIn2 = 32'd97; 
32'd693: dataIn2 = 32'd51; 
32'd694: dataIn2 = 32'd12; 
32'd695: dataIn2 = 32'd67; 
32'd696: dataIn2 = 32'd14; 
32'd697: dataIn2 = 32'd19; 
32'd698: dataIn2 = 32'd34; 
32'd699: dataIn2 = 32'd57; 
32'd700: dataIn2 = 32'd88; 
32'd701: dataIn2 = 32'd71; 
32'd702: dataIn2 = 32'd56; 
32'd703: dataIn2 = 32'd23; 
32'd704: dataIn2 = 32'd45; 
32'd705: dataIn2 = 32'd3; 
32'd706: dataIn2 = 32'd78; 
32'd707: dataIn2 = 32'd42; 
32'd708: dataIn2 = 32'd3; 
32'd709: dataIn2 = 32'd58; 
32'd710: dataIn2 = 32'd42; 
32'd711: dataIn2 = 32'd43; 
32'd712: dataIn2 = 32'd93; 
32'd713: dataIn2 = 32'd76; 
32'd714: dataIn2 = 32'd14; 
32'd715: dataIn2 = 32'd79; 
32'd716: dataIn2 = 32'd51; 
32'd717: dataIn2 = 32'd10; 
32'd718: dataIn2 = 32'd1; 
32'd719: dataIn2 = 32'd58; 
32'd720: dataIn2 = 32'd20; 
32'd721: dataIn2 = 32'd72; 
32'd722: dataIn2 = 32'd49; 
32'd723: dataIn2 = 32'd70; 
32'd724: dataIn2 = 32'd22; 
32'd725: dataIn2 = 32'd58; 
32'd726: dataIn2 = 32'd73; 
32'd727: dataIn2 = 32'd77; 
32'd728: dataIn2 = 32'd45; 
32'd729: dataIn2 = 32'd7; 
32'd730: dataIn2 = 32'd11; 
32'd731: dataIn2 = 32'd22; 
32'd732: dataIn2 = 32'd75; 
32'd733: dataIn2 = 32'd28; 
32'd734: dataIn2 = 32'd43; 
32'd735: dataIn2 = 32'd5; 
32'd736: dataIn2 = 32'd67; 
32'd737: dataIn2 = 32'd38; 
32'd738: dataIn2 = 32'd64; 
32'd739: dataIn2 = 32'd97; 
32'd740: dataIn2 = 32'd77; 
32'd741: dataIn2 = 32'd52; 
32'd742: dataIn2 = 32'd52; 
32'd743: dataIn2 = 32'd40; 
32'd744: dataIn2 = 32'd45; 
32'd745: dataIn2 = 32'd31; 
32'd746: dataIn2 = 32'd68; 
32'd747: dataIn2 = 32'd90; 
32'd748: dataIn2 = 32'd3; 
32'd749: dataIn2 = 32'd62; 
32'd750: dataIn2 = 32'd33; 
32'd751: dataIn2 = 32'd87; 
32'd752: dataIn2 = 32'd52; 
32'd753: dataIn2 = 32'd18; 
32'd754: dataIn2 = 32'd7; 
32'd755: dataIn2 = 32'd63; 
32'd756: dataIn2 = 32'd42; 
32'd757: dataIn2 = 32'd91; 
32'd758: dataIn2 = 32'd34; 
32'd759: dataIn2 = 32'd97; 
32'd760: dataIn2 = 32'd30; 
32'd761: dataIn2 = 32'd59; 
32'd762: dataIn2 = 32'd53; 
32'd763: dataIn2 = 32'd91; 
32'd764: dataIn2 = 32'd56; 
32'd765: dataIn2 = 32'd44; 
32'd766: dataIn2 = 32'd32; 
32'd767: dataIn2 = 32'd39; 
32'd768: dataIn2 = 32'd51; 
32'd769: dataIn2 = 32'd78; 
32'd770: dataIn2 = 32'd77; 
32'd771: dataIn2 = 32'd34; 
32'd772: dataIn2 = 32'd4; 
32'd773: dataIn2 = 32'd78; 
32'd774: dataIn2 = 32'd38; 
32'd775: dataIn2 = 32'd83; 
32'd776: dataIn2 = 32'd26; 
32'd777: dataIn2 = 32'd1; 
32'd778: dataIn2 = 32'd23; 
32'd779: dataIn2 = 32'd14; 
32'd780: dataIn2 = 32'd92; 
32'd781: dataIn2 = 32'd43; 
32'd782: dataIn2 = 32'd84; 
32'd783: dataIn2 = 32'd77; 
32'd784: dataIn2 = 32'd59; 
32'd785: dataIn2 = 32'd30; 
32'd786: dataIn2 = 32'd68; 
32'd787: dataIn2 = 32'd24; 
32'd788: dataIn2 = 32'd55; 
32'd789: dataIn2 = 32'd83; 
32'd790: dataIn2 = 32'd84; 
32'd791: dataIn2 = 32'd13; 
32'd792: dataIn2 = 32'd9; 
32'd793: dataIn2 = 32'd46; 
32'd794: dataIn2 = 32'd44; 
32'd795: dataIn2 = 32'd100; 
32'd796: dataIn2 = 32'd32; 
32'd797: dataIn2 = 32'd13; 
32'd798: dataIn2 = 32'd85; 
32'd799: dataIn2 = 32'd29; 
32'd800: dataIn2 = 32'd17; 
32'd801: dataIn2 = 32'd32; 
32'd802: dataIn2 = 32'd45; 
32'd803: dataIn2 = 32'd84; 
32'd804: dataIn2 = 32'd7; 
32'd805: dataIn2 = 32'd71; 
32'd806: dataIn2 = 32'd33; 
32'd807: dataIn2 = 32'd53; 
32'd808: dataIn2 = 32'd57; 
32'd809: dataIn2 = 32'd60; 
32'd810: dataIn2 = 32'd64; 
32'd811: dataIn2 = 32'd6; 
32'd812: dataIn2 = 32'd0; 
32'd813: dataIn2 = 32'd10; 
32'd814: dataIn2 = 32'd32; 
32'd815: dataIn2 = 32'd2; 
32'd816: dataIn2 = 32'd22; 
32'd817: dataIn2 = 32'd83; 
32'd818: dataIn2 = 32'd76; 
32'd819: dataIn2 = 32'd99; 
32'd820: dataIn2 = 32'd19; 
32'd821: dataIn2 = 32'd4; 
32'd822: dataIn2 = 32'd72; 
32'd823: dataIn2 = 32'd2; 
32'd824: dataIn2 = 32'd92; 
32'd825: dataIn2 = 32'd9; 
32'd826: dataIn2 = 32'd69; 
32'd827: dataIn2 = 32'd30; 
32'd828: dataIn2 = 32'd4; 
32'd829: dataIn2 = 32'd43; 
32'd830: dataIn2 = 32'd12; 
32'd831: dataIn2 = 32'd42; 
32'd832: dataIn2 = 32'd49; 
32'd833: dataIn2 = 32'd45; 
32'd834: dataIn2 = 32'd37; 
32'd835: dataIn2 = 32'd69; 
32'd836: dataIn2 = 32'd90; 
32'd837: dataIn2 = 32'd87; 
32'd838: dataIn2 = 32'd57; 
32'd839: dataIn2 = 32'd45; 
32'd840: dataIn2 = 32'd32; 
32'd841: dataIn2 = 32'd93; 
32'd842: dataIn2 = 32'd43; 
32'd843: dataIn2 = 32'd19; 
32'd844: dataIn2 = 32'd89; 
32'd845: dataIn2 = 32'd40; 
32'd846: dataIn2 = 32'd19; 
32'd847: dataIn2 = 32'd37; 
32'd848: dataIn2 = 32'd54; 
32'd849: dataIn2 = 32'd67; 
32'd850: dataIn2 = 32'd67; 
32'd851: dataIn2 = 32'd46; 
32'd852: dataIn2 = 32'd23; 
32'd853: dataIn2 = 32'd35; 
32'd854: dataIn2 = 32'd0; 
32'd855: dataIn2 = 32'd29; 
32'd856: dataIn2 = 32'd25; 
32'd857: dataIn2 = 32'd95; 
32'd858: dataIn2 = 32'd50; 
32'd859: dataIn2 = 32'd1; 
32'd860: dataIn2 = 32'd28; 
32'd861: dataIn2 = 32'd45; 
32'd862: dataIn2 = 32'd20; 
32'd863: dataIn2 = 32'd69; 
32'd864: dataIn2 = 32'd45; 
32'd865: dataIn2 = 32'd88; 
32'd866: dataIn2 = 32'd48; 
32'd867: dataIn2 = 32'd95; 
32'd868: dataIn2 = 32'd17; 
32'd869: dataIn2 = 32'd87; 
32'd870: dataIn2 = 32'd54; 
32'd871: dataIn2 = 32'd55; 
32'd872: dataIn2 = 32'd28; 
32'd873: dataIn2 = 32'd51; 
32'd874: dataIn2 = 32'd97; 
32'd875: dataIn2 = 32'd4; 
32'd876: dataIn2 = 32'd40; 
32'd877: dataIn2 = 32'd67; 
32'd878: dataIn2 = 32'd92; 
32'd879: dataIn2 = 32'd42; 
32'd880: dataIn2 = 32'd79; 
32'd881: dataIn2 = 32'd63; 
32'd882: dataIn2 = 32'd18; 
32'd883: dataIn2 = 32'd5; 
32'd884: dataIn2 = 32'd77; 
32'd885: dataIn2 = 32'd82; 
32'd886: dataIn2 = 32'd27; 
32'd887: dataIn2 = 32'd74; 
32'd888: dataIn2 = 32'd83; 
32'd889: dataIn2 = 32'd44; 
32'd890: dataIn2 = 32'd5; 
32'd891: dataIn2 = 32'd42; 
32'd892: dataIn2 = 32'd11; 
32'd893: dataIn2 = 32'd89; 
32'd894: dataIn2 = 32'd70; 
32'd895: dataIn2 = 32'd44; 
32'd896: dataIn2 = 32'd7; 
32'd897: dataIn2 = 32'd75; 
32'd898: dataIn2 = 32'd66; 
32'd899: dataIn2 = 32'd79; 
32'd900: dataIn2 = 32'd36; 
32'd901: dataIn2 = 32'd71; 
32'd902: dataIn2 = 32'd66; 
32'd903: dataIn2 = 32'd80; 
32'd904: dataIn2 = 32'd89; 
32'd905: dataIn2 = 32'd92; 
32'd906: dataIn2 = 32'd3; 
32'd907: dataIn2 = 32'd33; 
32'd908: dataIn2 = 32'd99; 
32'd909: dataIn2 = 32'd15; 
32'd910: dataIn2 = 32'd74; 
32'd911: dataIn2 = 32'd44; 
32'd912: dataIn2 = 32'd53; 
32'd913: dataIn2 = 32'd86; 
32'd914: dataIn2 = 32'd50; 
32'd915: dataIn2 = 32'd5; 
32'd916: dataIn2 = 32'd1; 
32'd917: dataIn2 = 32'd51; 
32'd918: dataIn2 = 32'd76; 
32'd919: dataIn2 = 32'd32; 
32'd920: dataIn2 = 32'd59; 
32'd921: dataIn2 = 32'd21; 
32'd922: dataIn2 = 32'd15; 
32'd923: dataIn2 = 32'd79; 
32'd924: dataIn2 = 32'd96; 
32'd925: dataIn2 = 32'd51; 
32'd926: dataIn2 = 32'd6; 
32'd927: dataIn2 = 32'd68; 
32'd928: dataIn2 = 32'd13; 
32'd929: dataIn2 = 32'd97; 
32'd930: dataIn2 = 32'd36; 
32'd931: dataIn2 = 32'd82; 
32'd932: dataIn2 = 32'd23; 
32'd933: dataIn2 = 32'd91; 
32'd934: dataIn2 = 32'd79; 
32'd935: dataIn2 = 32'd12; 
32'd936: dataIn2 = 32'd59; 
32'd937: dataIn2 = 32'd28; 
32'd938: dataIn2 = 32'd22; 
32'd939: dataIn2 = 32'd85; 
32'd940: dataIn2 = 32'd77; 
32'd941: dataIn2 = 32'd16; 
32'd942: dataIn2 = 32'd86; 
32'd943: dataIn2 = 32'd66; 
32'd944: dataIn2 = 32'd55; 
32'd945: dataIn2 = 32'd43; 
32'd946: dataIn2 = 32'd25; 
32'd947: dataIn2 = 32'd72; 
32'd948: dataIn2 = 32'd93; 
32'd949: dataIn2 = 32'd67; 
32'd950: dataIn2 = 32'd45; 
32'd951: dataIn2 = 32'd69; 
32'd952: dataIn2 = 32'd48; 
32'd953: dataIn2 = 32'd78; 
32'd954: dataIn2 = 32'd16; 
32'd955: dataIn2 = 32'd52; 
32'd956: dataIn2 = 32'd7; 
32'd957: dataIn2 = 32'd61; 
32'd958: dataIn2 = 32'd51; 
32'd959: dataIn2 = 32'd55; 
32'd960: dataIn2 = 32'd17; 
32'd961: dataIn2 = 32'd82; 
32'd962: dataIn2 = 32'd38; 
32'd963: dataIn2 = 32'd52; 
32'd964: dataIn2 = 32'd99; 
32'd965: dataIn2 = 32'd77; 
32'd966: dataIn2 = 32'd23; 
32'd967: dataIn2 = 32'd78; 
32'd968: dataIn2 = 32'd32; 
32'd969: dataIn2 = 32'd45; 
32'd970: dataIn2 = 32'd94; 
32'd971: dataIn2 = 32'd97; 
32'd972: dataIn2 = 32'd87; 
32'd973: dataIn2 = 32'd2; 
32'd974: dataIn2 = 32'd49; 
32'd975: dataIn2 = 32'd92; 
32'd976: dataIn2 = 32'd41; 
32'd977: dataIn2 = 32'd77; 
32'd978: dataIn2 = 32'd35; 
32'd979: dataIn2 = 32'd45; 
32'd980: dataIn2 = 32'd87; 
32'd981: dataIn2 = 32'd26; 
32'd982: dataIn2 = 32'd96; 
32'd983: dataIn2 = 32'd66; 
32'd984: dataIn2 = 32'd1; 
32'd985: dataIn2 = 32'd19; 
32'd986: dataIn2 = 32'd77; 
32'd987: dataIn2 = 32'd73; 
32'd988: dataIn2 = 32'd27; 
32'd989: dataIn2 = 32'd40; 
32'd990: dataIn2 = 32'd43; 
32'd991: dataIn2 = 32'd50; 
32'd992: dataIn2 = 32'd82; 
32'd993: dataIn2 = 32'd10; 
32'd994: dataIn2 = 32'd33; 
32'd995: dataIn2 = 32'd71; 
32'd996: dataIn2 = 32'd63; 
32'd997: dataIn2 = 32'd5; 
32'd998: dataIn2 = 32'd27; 
32'd999: dataIn2 = 32'd34; 
32'd1000: dataIn2 = 32'd81; 
32'd1001: dataIn2 = 32'd71; 
32'd1002: dataIn2 = 32'd87; 
32'd1003: dataIn2 = 32'd99; 
32'd1004: dataIn2 = 32'd16; 
32'd1005: dataIn2 = 32'd70; 
32'd1006: dataIn2 = 32'd81; 
32'd1007: dataIn2 = 32'd18; 
32'd1008: dataIn2 = 32'd67; 
32'd1009: dataIn2 = 32'd36; 
32'd1010: dataIn2 = 32'd15; 
32'd1011: dataIn2 = 32'd84; 
32'd1012: dataIn2 = 32'd76; 
32'd1013: dataIn2 = 32'd8; 
32'd1014: dataIn2 = 32'd64; 
32'd1015: dataIn2 = 32'd66; 
32'd1016: dataIn2 = 32'd95; 
32'd1017: dataIn2 = 32'd92; 
32'd1018: dataIn2 = 32'd99; 
32'd1019: dataIn2 = 32'd77; 
32'd1020: dataIn2 = 32'd41; 
32'd1021: dataIn2 = 32'd24; 
32'd1022: dataIn2 = 32'd84; 
32'd1023: dataIn2 = 32'd46; 
32'd1024: dataIn2 = 32'd36; 
32'd1025: dataIn2 = 32'd73; 
32'd1026: dataIn2 = 32'd45; 
32'd1027: dataIn2 = 32'd93; 
32'd1028: dataIn2 = 32'd76; 
32'd1029: dataIn2 = 32'd45; 
32'd1030: dataIn2 = 32'd55; 
32'd1031: dataIn2 = 32'd68; 
32'd1032: dataIn2 = 32'd31; 
32'd1033: dataIn2 = 32'd2; 
32'd1034: dataIn2 = 32'd98; 
32'd1035: dataIn2 = 32'd14; 
32'd1036: dataIn2 = 32'd17; 
32'd1037: dataIn2 = 32'd62; 
32'd1038: dataIn2 = 32'd99; 
32'd1039: dataIn2 = 32'd94; 
32'd1040: dataIn2 = 32'd86; 
32'd1041: dataIn2 = 32'd7; 
32'd1042: dataIn2 = 32'd61; 
32'd1043: dataIn2 = 32'd46; 
32'd1044: dataIn2 = 32'd41; 
32'd1045: dataIn2 = 32'd19; 
32'd1046: dataIn2 = 32'd19; 
32'd1047: dataIn2 = 32'd5; 
32'd1048: dataIn2 = 32'd56; 
32'd1049: dataIn2 = 32'd82; 
32'd1050: dataIn2 = 32'd23; 
32'd1051: dataIn2 = 32'd95; 
32'd1052: dataIn2 = 32'd97; 
32'd1053: dataIn2 = 32'd94; 
32'd1054: dataIn2 = 32'd41; 
32'd1055: dataIn2 = 32'd25; 
32'd1056: dataIn2 = 32'd52; 
32'd1057: dataIn2 = 32'd55; 
32'd1058: dataIn2 = 32'd87; 
32'd1059: dataIn2 = 32'd30; 
32'd1060: dataIn2 = 32'd45; 
32'd1061: dataIn2 = 32'd18; 
32'd1062: dataIn2 = 32'd78; 
32'd1063: dataIn2 = 32'd99; 
32'd1064: dataIn2 = 32'd92; 
32'd1065: dataIn2 = 32'd90; 
32'd1066: dataIn2 = 32'd31; 
32'd1067: dataIn2 = 32'd5; 
32'd1068: dataIn2 = 32'd12; 
32'd1069: dataIn2 = 32'd47; 
32'd1070: dataIn2 = 32'd82; 
32'd1071: dataIn2 = 32'd14; 
32'd1072: dataIn2 = 32'd58; 
32'd1073: dataIn2 = 32'd96; 
32'd1074: dataIn2 = 32'd88; 
32'd1075: dataIn2 = 32'd59; 
32'd1076: dataIn2 = 32'd69; 
32'd1077: dataIn2 = 32'd58; 
32'd1078: dataIn2 = 32'd44; 
32'd1079: dataIn2 = 32'd33; 
32'd1080: dataIn2 = 32'd87; 
32'd1081: dataIn2 = 32'd94; 
32'd1082: dataIn2 = 32'd53; 
32'd1083: dataIn2 = 32'd31; 
32'd1084: dataIn2 = 32'd86; 
32'd1085: dataIn2 = 32'd28; 
32'd1086: dataIn2 = 32'd28; 
32'd1087: dataIn2 = 32'd85; 
32'd1088: dataIn2 = 32'd59; 
32'd1089: dataIn2 = 32'd33; 
32'd1090: dataIn2 = 32'd3; 
32'd1091: dataIn2 = 32'd77; 
32'd1092: dataIn2 = 32'd52; 
32'd1093: dataIn2 = 32'd92; 
32'd1094: dataIn2 = 32'd56; 
32'd1095: dataIn2 = 32'd96; 
32'd1096: dataIn2 = 32'd22; 
32'd1097: dataIn2 = 32'd0; 
32'd1098: dataIn2 = 32'd4; 
32'd1099: dataIn2 = 32'd2; 
32'd1100: dataIn2 = 32'd44; 
32'd1101: dataIn2 = 32'd31; 
32'd1102: dataIn2 = 32'd60; 
32'd1103: dataIn2 = 32'd43; 
32'd1104: dataIn2 = 32'd68; 
32'd1105: dataIn2 = 32'd47; 
32'd1106: dataIn2 = 32'd14; 
32'd1107: dataIn2 = 32'd75; 
32'd1108: dataIn2 = 32'd40; 
32'd1109: dataIn2 = 32'd51; 
32'd1110: dataIn2 = 32'd12; 
32'd1111: dataIn2 = 32'd79; 
32'd1112: dataIn2 = 32'd71; 
32'd1113: dataIn2 = 32'd73; 
32'd1114: dataIn2 = 32'd56; 
32'd1115: dataIn2 = 32'd63; 
32'd1116: dataIn2 = 32'd88; 
32'd1117: dataIn2 = 32'd4; 
32'd1118: dataIn2 = 32'd78; 
32'd1119: dataIn2 = 32'd75; 
32'd1120: dataIn2 = 32'd51; 
32'd1121: dataIn2 = 32'd63; 
32'd1122: dataIn2 = 32'd59; 
32'd1123: dataIn2 = 32'd90; 
32'd1124: dataIn2 = 32'd53; 
32'd1125: dataIn2 = 32'd11; 
32'd1126: dataIn2 = 32'd51; 
32'd1127: dataIn2 = 32'd83; 
32'd1128: dataIn2 = 32'd80; 
32'd1129: dataIn2 = 32'd59; 
32'd1130: dataIn2 = 32'd53; 
32'd1131: dataIn2 = 32'd4; 
32'd1132: dataIn2 = 32'd39; 
32'd1133: dataIn2 = 32'd27; 
32'd1134: dataIn2 = 32'd12; 
32'd1135: dataIn2 = 32'd76; 
32'd1136: dataIn2 = 32'd52; 
32'd1137: dataIn2 = 32'd43; 
32'd1138: dataIn2 = 32'd74; 
32'd1139: dataIn2 = 32'd72; 
32'd1140: dataIn2 = 32'd7; 
32'd1141: dataIn2 = 32'd45; 
32'd1142: dataIn2 = 32'd46; 
32'd1143: dataIn2 = 32'd54; 
32'd1144: dataIn2 = 32'd44; 
32'd1145: dataIn2 = 32'd13; 
32'd1146: dataIn2 = 32'd35; 
32'd1147: dataIn2 = 32'd4; 
32'd1148: dataIn2 = 32'd79; 
32'd1149: dataIn2 = 32'd92; 
32'd1150: dataIn2 = 32'd15; 
32'd1151: dataIn2 = 32'd10; 
32'd1152: dataIn2 = 32'd74; 
32'd1153: dataIn2 = 32'd77; 
32'd1154: dataIn2 = 32'd86; 
32'd1155: dataIn2 = 32'd64; 
32'd1156: dataIn2 = 32'd2; 
32'd1157: dataIn2 = 32'd90; 
32'd1158: dataIn2 = 32'd78; 
32'd1159: dataIn2 = 32'd5; 
32'd1160: dataIn2 = 32'd6; 
32'd1161: dataIn2 = 32'd38; 
32'd1162: dataIn2 = 32'd10; 
32'd1163: dataIn2 = 32'd82; 
32'd1164: dataIn2 = 32'd35; 
32'd1165: dataIn2 = 32'd71; 
32'd1166: dataIn2 = 32'd64; 
32'd1167: dataIn2 = 32'd5; 
32'd1168: dataIn2 = 32'd50; 
32'd1169: dataIn2 = 32'd10; 
32'd1170: dataIn2 = 32'd59; 
32'd1171: dataIn2 = 32'd23; 
32'd1172: dataIn2 = 32'd33; 
32'd1173: dataIn2 = 32'd81; 
32'd1174: dataIn2 = 32'd13; 
32'd1175: dataIn2 = 32'd64; 
32'd1176: dataIn2 = 32'd23; 
32'd1177: dataIn2 = 32'd29; 
32'd1178: dataIn2 = 32'd54; 
32'd1179: dataIn2 = 32'd39; 
32'd1180: dataIn2 = 32'd49; 
32'd1181: dataIn2 = 32'd72; 
32'd1182: dataIn2 = 32'd63; 
32'd1183: dataIn2 = 32'd99; 
32'd1184: dataIn2 = 32'd72; 
32'd1185: dataIn2 = 32'd48; 
32'd1186: dataIn2 = 32'd36; 
32'd1187: dataIn2 = 32'd51; 
32'd1188: dataIn2 = 32'd26; 
32'd1189: dataIn2 = 32'd14; 
32'd1190: dataIn2 = 32'd94; 
32'd1191: dataIn2 = 32'd69; 
32'd1192: dataIn2 = 32'd67; 
32'd1193: dataIn2 = 32'd14; 
32'd1194: dataIn2 = 32'd93; 
32'd1195: dataIn2 = 32'd37; 
32'd1196: dataIn2 = 32'd94; 
32'd1197: dataIn2 = 32'd11; 
32'd1198: dataIn2 = 32'd24; 
32'd1199: dataIn2 = 32'd21; 
32'd1200: dataIn2 = 32'd25; 
32'd1201: dataIn2 = 32'd95; 
32'd1202: dataIn2 = 32'd4; 
32'd1203: dataIn2 = 32'd73; 
32'd1204: dataIn2 = 32'd85; 
32'd1205: dataIn2 = 32'd68; 
32'd1206: dataIn2 = 32'd58; 
32'd1207: dataIn2 = 32'd29; 
32'd1208: dataIn2 = 32'd74; 
32'd1209: dataIn2 = 32'd20; 
32'd1210: dataIn2 = 32'd72; 
32'd1211: dataIn2 = 32'd100; 
32'd1212: dataIn2 = 32'd84; 
32'd1213: dataIn2 = 32'd71; 
32'd1214: dataIn2 = 32'd5; 
32'd1215: dataIn2 = 32'd34; 
32'd1216: dataIn2 = 32'd22; 
32'd1217: dataIn2 = 32'd32; 
32'd1218: dataIn2 = 32'd35; 
32'd1219: dataIn2 = 32'd2; 
32'd1220: dataIn2 = 32'd55; 
32'd1221: dataIn2 = 32'd39; 
32'd1222: dataIn2 = 32'd58; 
32'd1223: dataIn2 = 32'd73; 
32'd1224: dataIn2 = 32'd30; 
32'd1225: dataIn2 = 32'd58; 
32'd1226: dataIn2 = 32'd9; 
32'd1227: dataIn2 = 32'd29; 
32'd1228: dataIn2 = 32'd96; 
32'd1229: dataIn2 = 32'd9; 
32'd1230: dataIn2 = 32'd82; 
32'd1231: dataIn2 = 32'd19; 
32'd1232: dataIn2 = 32'd59; 
32'd1233: dataIn2 = 32'd36; 
32'd1234: dataIn2 = 32'd21; 
32'd1235: dataIn2 = 32'd7; 
32'd1236: dataIn2 = 32'd70; 
32'd1237: dataIn2 = 32'd8; 
32'd1238: dataIn2 = 32'd56; 
32'd1239: dataIn2 = 32'd5; 
32'd1240: dataIn2 = 32'd28; 
32'd1241: dataIn2 = 32'd69; 
32'd1242: dataIn2 = 32'd93; 
32'd1243: dataIn2 = 32'd60; 
32'd1244: dataIn2 = 32'd0; 
32'd1245: dataIn2 = 32'd82; 
32'd1246: dataIn2 = 32'd90; 
32'd1247: dataIn2 = 32'd39; 
32'd1248: dataIn2 = 32'd78; 
32'd1249: dataIn2 = 32'd95; 
32'd1250: dataIn2 = 32'd76; 
32'd1251: dataIn2 = 32'd19; 
32'd1252: dataIn2 = 32'd16; 
32'd1253: dataIn2 = 32'd22; 
32'd1254: dataIn2 = 32'd99; 
32'd1255: dataIn2 = 32'd74; 
32'd1256: dataIn2 = 32'd50; 
32'd1257: dataIn2 = 32'd95; 
32'd1258: dataIn2 = 32'd70; 
32'd1259: dataIn2 = 32'd58; 
32'd1260: dataIn2 = 32'd53; 
32'd1261: dataIn2 = 32'd100; 
32'd1262: dataIn2 = 32'd60; 
32'd1263: dataIn2 = 32'd29; 
32'd1264: dataIn2 = 32'd71; 
32'd1265: dataIn2 = 32'd40; 
32'd1266: dataIn2 = 32'd40; 
32'd1267: dataIn2 = 32'd44; 
32'd1268: dataIn2 = 32'd87; 
32'd1269: dataIn2 = 32'd72; 
32'd1270: dataIn2 = 32'd46; 
32'd1271: dataIn2 = 32'd14; 
32'd1272: dataIn2 = 32'd22; 
32'd1273: dataIn2 = 32'd18; 
32'd1274: dataIn2 = 32'd33; 
32'd1275: dataIn2 = 32'd50; 
32'd1276: dataIn2 = 32'd9; 
32'd1277: dataIn2 = 32'd91; 
32'd1278: dataIn2 = 32'd11; 
32'd1279: dataIn2 = 32'd97; 
32'd1280: dataIn2 = 32'd75; 
32'd1281: dataIn2 = 32'd77; 
32'd1282: dataIn2 = 32'd63; 
32'd1283: dataIn2 = 32'd38; 
32'd1284: dataIn2 = 32'd69; 
32'd1285: dataIn2 = 32'd43; 
32'd1286: dataIn2 = 32'd52; 
32'd1287: dataIn2 = 32'd41; 
32'd1288: dataIn2 = 32'd35; 
32'd1289: dataIn2 = 32'd52; 
32'd1290: dataIn2 = 32'd71; 
32'd1291: dataIn2 = 32'd67; 
32'd1292: dataIn2 = 32'd22; 
32'd1293: dataIn2 = 32'd49; 
32'd1294: dataIn2 = 32'd27; 
32'd1295: dataIn2 = 32'd72; 
32'd1296: dataIn2 = 32'd26; 
32'd1297: dataIn2 = 32'd94; 
32'd1298: dataIn2 = 32'd40; 
32'd1299: dataIn2 = 32'd63; 
32'd1300: dataIn2 = 32'd73; 
32'd1301: dataIn2 = 32'd82; 
32'd1302: dataIn2 = 32'd69; 
32'd1303: dataIn2 = 32'd53; 
32'd1304: dataIn2 = 32'd44; 
32'd1305: dataIn2 = 32'd0; 
32'd1306: dataIn2 = 32'd51; 
32'd1307: dataIn2 = 32'd82; 
32'd1308: dataIn2 = 32'd51; 
32'd1309: dataIn2 = 32'd79; 
32'd1310: dataIn2 = 32'd5; 
32'd1311: dataIn2 = 32'd10; 
32'd1312: dataIn2 = 32'd5; 
32'd1313: dataIn2 = 32'd16; 
32'd1314: dataIn2 = 32'd39; 
32'd1315: dataIn2 = 32'd50; 
32'd1316: dataIn2 = 32'd70; 
32'd1317: dataIn2 = 32'd30; 
32'd1318: dataIn2 = 32'd31; 
32'd1319: dataIn2 = 32'd92; 
32'd1320: dataIn2 = 32'd32; 
32'd1321: dataIn2 = 32'd44; 
32'd1322: dataIn2 = 32'd4; 
32'd1323: dataIn2 = 32'd33; 
32'd1324: dataIn2 = 32'd33; 
32'd1325: dataIn2 = 32'd97; 
32'd1326: dataIn2 = 32'd85; 
32'd1327: dataIn2 = 32'd34; 
32'd1328: dataIn2 = 32'd11; 
32'd1329: dataIn2 = 32'd24; 
32'd1330: dataIn2 = 32'd75; 
32'd1331: dataIn2 = 32'd37; 
32'd1332: dataIn2 = 32'd62; 
32'd1333: dataIn2 = 32'd100; 
32'd1334: dataIn2 = 32'd79; 
32'd1335: dataIn2 = 32'd25; 
32'd1336: dataIn2 = 32'd5; 
32'd1337: dataIn2 = 32'd45; 
32'd1338: dataIn2 = 32'd94; 
32'd1339: dataIn2 = 32'd55; 
32'd1340: dataIn2 = 32'd7; 
32'd1341: dataIn2 = 32'd85; 
32'd1342: dataIn2 = 32'd79; 
32'd1343: dataIn2 = 32'd26; 
32'd1344: dataIn2 = 32'd2; 
32'd1345: dataIn2 = 32'd17; 
32'd1346: dataIn2 = 32'd93; 
32'd1347: dataIn2 = 32'd98; 
32'd1348: dataIn2 = 32'd57; 
32'd1349: dataIn2 = 32'd21; 
32'd1350: dataIn2 = 32'd87; 
32'd1351: dataIn2 = 32'd61; 
32'd1352: dataIn2 = 32'd1; 
32'd1353: dataIn2 = 32'd11; 
32'd1354: dataIn2 = 32'd64; 
32'd1355: dataIn2 = 32'd29; 
32'd1356: dataIn2 = 32'd26; 
32'd1357: dataIn2 = 32'd96; 
32'd1358: dataIn2 = 32'd61; 
32'd1359: dataIn2 = 32'd44; 
32'd1360: dataIn2 = 32'd49; 
32'd1361: dataIn2 = 32'd4; 
32'd1362: dataIn2 = 32'd44; 
32'd1363: dataIn2 = 32'd24; 
32'd1364: dataIn2 = 32'd3; 
32'd1365: dataIn2 = 32'd26; 
32'd1366: dataIn2 = 32'd92; 
32'd1367: dataIn2 = 32'd53; 
32'd1368: dataIn2 = 32'd43; 
32'd1369: dataIn2 = 32'd54; 
32'd1370: dataIn2 = 32'd81; 
32'd1371: dataIn2 = 32'd13; 
32'd1372: dataIn2 = 32'd18; 
32'd1373: dataIn2 = 32'd18; 
32'd1374: dataIn2 = 32'd76; 
32'd1375: dataIn2 = 32'd93; 
32'd1376: dataIn2 = 32'd53; 
32'd1377: dataIn2 = 32'd66; 
32'd1378: dataIn2 = 32'd39; 
32'd1379: dataIn2 = 32'd51; 
32'd1380: dataIn2 = 32'd29; 
32'd1381: dataIn2 = 32'd29; 
32'd1382: dataIn2 = 32'd3; 
32'd1383: dataIn2 = 32'd90; 
32'd1384: dataIn2 = 32'd73; 
32'd1385: dataIn2 = 32'd49; 
32'd1386: dataIn2 = 32'd4; 
32'd1387: dataIn2 = 32'd66; 
32'd1388: dataIn2 = 32'd74; 
32'd1389: dataIn2 = 32'd69; 
32'd1390: dataIn2 = 32'd11; 
32'd1391: dataIn2 = 32'd71; 
32'd1392: dataIn2 = 32'd42; 
32'd1393: dataIn2 = 32'd39; 
32'd1394: dataIn2 = 32'd100; 
32'd1395: dataIn2 = 32'd58; 
32'd1396: dataIn2 = 32'd68; 
32'd1397: dataIn2 = 32'd18; 
32'd1398: dataIn2 = 32'd22; 
32'd1399: dataIn2 = 32'd16; 
32'd1400: dataIn2 = 32'd22; 
32'd1401: dataIn2 = 32'd6; 
32'd1402: dataIn2 = 32'd66; 
32'd1403: dataIn2 = 32'd18; 
32'd1404: dataIn2 = 32'd31; 
32'd1405: dataIn2 = 32'd78; 
32'd1406: dataIn2 = 32'd71; 
32'd1407: dataIn2 = 32'd90; 
32'd1408: dataIn2 = 32'd78; 
32'd1409: dataIn2 = 32'd34; 
32'd1410: dataIn2 = 32'd36; 
32'd1411: dataIn2 = 32'd60; 
32'd1412: dataIn2 = 32'd47; 
32'd1413: dataIn2 = 32'd39; 
32'd1414: dataIn2 = 32'd29; 
32'd1415: dataIn2 = 32'd89; 
32'd1416: dataIn2 = 32'd99; 
32'd1417: dataIn2 = 32'd74; 
32'd1418: dataIn2 = 32'd16; 
32'd1419: dataIn2 = 32'd54; 
32'd1420: dataIn2 = 32'd100; 
32'd1421: dataIn2 = 32'd65; 
32'd1422: dataIn2 = 32'd6; 
32'd1423: dataIn2 = 32'd65; 
32'd1424: dataIn2 = 32'd83; 
32'd1425: dataIn2 = 32'd24; 
32'd1426: dataIn2 = 32'd32; 
32'd1427: dataIn2 = 32'd95; 
32'd1428: dataIn2 = 32'd73; 
32'd1429: dataIn2 = 32'd58; 
32'd1430: dataIn2 = 32'd71; 
32'd1431: dataIn2 = 32'd1; 
32'd1432: dataIn2 = 32'd30; 
32'd1433: dataIn2 = 32'd36; 
32'd1434: dataIn2 = 32'd92; 
32'd1435: dataIn2 = 32'd67; 
32'd1436: dataIn2 = 32'd85; 
32'd1437: dataIn2 = 32'd56; 
32'd1438: dataIn2 = 32'd4; 
32'd1439: dataIn2 = 32'd60; 
32'd1440: dataIn2 = 32'd87; 
32'd1441: dataIn2 = 32'd8; 
32'd1442: dataIn2 = 32'd54; 
32'd1443: dataIn2 = 32'd11; 
32'd1444: dataIn2 = 32'd1; 
32'd1445: dataIn2 = 32'd30; 
32'd1446: dataIn2 = 32'd8; 
32'd1447: dataIn2 = 32'd81; 
32'd1448: dataIn2 = 32'd11; 
32'd1449: dataIn2 = 32'd41; 
32'd1450: dataIn2 = 32'd70; 
32'd1451: dataIn2 = 32'd45; 
32'd1452: dataIn2 = 32'd73; 
32'd1453: dataIn2 = 32'd98; 
32'd1454: dataIn2 = 32'd29; 
32'd1455: dataIn2 = 32'd83; 
32'd1456: dataIn2 = 32'd55; 
32'd1457: dataIn2 = 32'd96; 
32'd1458: dataIn2 = 32'd81; 
32'd1459: dataIn2 = 32'd11; 
32'd1460: dataIn2 = 32'd57; 
32'd1461: dataIn2 = 32'd51; 
32'd1462: dataIn2 = 32'd26; 
32'd1463: dataIn2 = 32'd5; 
32'd1464: dataIn2 = 32'd70; 
32'd1465: dataIn2 = 32'd72; 
32'd1466: dataIn2 = 32'd55; 
32'd1467: dataIn2 = 32'd62; 
32'd1468: dataIn2 = 32'd61; 
32'd1469: dataIn2 = 32'd33; 
32'd1470: dataIn2 = 32'd80; 
32'd1471: dataIn2 = 32'd99; 
32'd1472: dataIn2 = 32'd46; 
32'd1473: dataIn2 = 32'd82; 
32'd1474: dataIn2 = 32'd29; 
32'd1475: dataIn2 = 32'd89; 
32'd1476: dataIn2 = 32'd93; 
32'd1477: dataIn2 = 32'd6; 
32'd1478: dataIn2 = 32'd78; 
32'd1479: dataIn2 = 32'd34; 
32'd1480: dataIn2 = 32'd34; 
32'd1481: dataIn2 = 32'd70; 
32'd1482: dataIn2 = 32'd81; 
32'd1483: dataIn2 = 32'd31; 
32'd1484: dataIn2 = 32'd43; 
32'd1485: dataIn2 = 32'd22; 
32'd1486: dataIn2 = 32'd89; 
32'd1487: dataIn2 = 32'd24; 
32'd1488: dataIn2 = 32'd50; 
32'd1489: dataIn2 = 32'd38; 
32'd1490: dataIn2 = 32'd72; 
32'd1491: dataIn2 = 32'd34; 
32'd1492: dataIn2 = 32'd63; 
32'd1493: dataIn2 = 32'd69; 
32'd1494: dataIn2 = 32'd14; 
32'd1495: dataIn2 = 32'd54; 
32'd1496: dataIn2 = 32'd44; 
32'd1497: dataIn2 = 32'd5; 
32'd1498: dataIn2 = 32'd92; 
32'd1499: dataIn2 = 32'd70; 
32'd1500: dataIn2 = 32'd6; 
32'd1501: dataIn2 = 32'd79; 
32'd1502: dataIn2 = 32'd56; 
32'd1503: dataIn2 = 32'd33; 
32'd1504: dataIn2 = 32'd2; 
32'd1505: dataIn2 = 32'd48; 
32'd1506: dataIn2 = 32'd39; 
32'd1507: dataIn2 = 32'd76; 
32'd1508: dataIn2 = 32'd95; 
32'd1509: dataIn2 = 32'd97; 
32'd1510: dataIn2 = 32'd12; 
32'd1511: dataIn2 = 32'd49; 
32'd1512: dataIn2 = 32'd7; 
32'd1513: dataIn2 = 32'd44; 
32'd1514: dataIn2 = 32'd51; 
32'd1515: dataIn2 = 32'd60; 
32'd1516: dataIn2 = 32'd89; 
32'd1517: dataIn2 = 32'd59; 
32'd1518: dataIn2 = 32'd0; 
32'd1519: dataIn2 = 32'd29; 
32'd1520: dataIn2 = 32'd11; 
32'd1521: dataIn2 = 32'd76; 
32'd1522: dataIn2 = 32'd79; 
32'd1523: dataIn2 = 32'd70; 
32'd1524: dataIn2 = 32'd3; 
32'd1525: dataIn2 = 32'd72; 
32'd1526: dataIn2 = 32'd53; 
32'd1527: dataIn2 = 32'd64; 
32'd1528: dataIn2 = 32'd55; 
32'd1529: dataIn2 = 32'd26; 
32'd1530: dataIn2 = 32'd49; 
32'd1531: dataIn2 = 32'd35; 
32'd1532: dataIn2 = 32'd62; 
32'd1533: dataIn2 = 32'd85; 
32'd1534: dataIn2 = 32'd42; 
32'd1535: dataIn2 = 32'd51; 
32'd1536: dataIn2 = 32'd66; 
32'd1537: dataIn2 = 32'd51; 
32'd1538: dataIn2 = 32'd65; 
32'd1539: dataIn2 = 32'd76; 
32'd1540: dataIn2 = 32'd63; 
32'd1541: dataIn2 = 32'd4; 
32'd1542: dataIn2 = 32'd12; 
32'd1543: dataIn2 = 32'd29; 
32'd1544: dataIn2 = 32'd55; 
32'd1545: dataIn2 = 32'd27; 
32'd1546: dataIn2 = 32'd41; 
32'd1547: dataIn2 = 32'd88; 
32'd1548: dataIn2 = 32'd89; 
32'd1549: dataIn2 = 32'd59; 
32'd1550: dataIn2 = 32'd82; 
32'd1551: dataIn2 = 32'd23; 
32'd1552: dataIn2 = 32'd33; 
32'd1553: dataIn2 = 32'd60; 
32'd1554: dataIn2 = 32'd50; 
32'd1555: dataIn2 = 32'd32; 
32'd1556: dataIn2 = 32'd19; 
32'd1557: dataIn2 = 32'd30; 
32'd1558: dataIn2 = 32'd25; 
32'd1559: dataIn2 = 32'd90; 
32'd1560: dataIn2 = 32'd9; 
32'd1561: dataIn2 = 32'd61; 
32'd1562: dataIn2 = 32'd28; 
32'd1563: dataIn2 = 32'd47; 
32'd1564: dataIn2 = 32'd48; 
32'd1565: dataIn2 = 32'd96; 
32'd1566: dataIn2 = 32'd60; 
32'd1567: dataIn2 = 32'd24; 
32'd1568: dataIn2 = 32'd96; 
32'd1569: dataIn2 = 32'd17; 
32'd1570: dataIn2 = 32'd13; 
32'd1571: dataIn2 = 32'd85; 
32'd1572: dataIn2 = 32'd30; 
32'd1573: dataIn2 = 32'd38; 
32'd1574: dataIn2 = 32'd18; 
32'd1575: dataIn2 = 32'd32; 
32'd1576: dataIn2 = 32'd63; 
32'd1577: dataIn2 = 32'd28; 
32'd1578: dataIn2 = 32'd78; 
32'd1579: dataIn2 = 32'd59; 
32'd1580: dataIn2 = 32'd62; 
32'd1581: dataIn2 = 32'd98; 
32'd1582: dataIn2 = 32'd91; 
32'd1583: dataIn2 = 32'd95; 
32'd1584: dataIn2 = 32'd67; 
32'd1585: dataIn2 = 32'd62; 
32'd1586: dataIn2 = 32'd26; 
32'd1587: dataIn2 = 32'd66; 
32'd1588: dataIn2 = 32'd25; 
32'd1589: dataIn2 = 32'd49; 
32'd1590: dataIn2 = 32'd88; 
32'd1591: dataIn2 = 32'd23; 
32'd1592: dataIn2 = 32'd3; 
32'd1593: dataIn2 = 32'd45; 
32'd1594: dataIn2 = 32'd13; 
32'd1595: dataIn2 = 32'd6; 
32'd1596: dataIn2 = 32'd99; 
32'd1597: dataIn2 = 32'd46; 
32'd1598: dataIn2 = 32'd34; 
32'd1599: dataIn2 = 32'd37; 
32'd1600: dataIn2 = 32'd87; 
32'd1601: dataIn2 = 32'd55; 
32'd1602: dataIn2 = 32'd45; 
32'd1603: dataIn2 = 32'd3; 
32'd1604: dataIn2 = 32'd38; 
32'd1605: dataIn2 = 32'd13; 
32'd1606: dataIn2 = 32'd64; 
32'd1607: dataIn2 = 32'd88; 
32'd1608: dataIn2 = 32'd10; 
32'd1609: dataIn2 = 32'd11; 
32'd1610: dataIn2 = 32'd52; 
32'd1611: dataIn2 = 32'd41; 
32'd1612: dataIn2 = 32'd12; 
32'd1613: dataIn2 = 32'd36; 
32'd1614: dataIn2 = 32'd65; 
32'd1615: dataIn2 = 32'd39; 
32'd1616: dataIn2 = 32'd46; 
32'd1617: dataIn2 = 32'd19; 
32'd1618: dataIn2 = 32'd71; 
32'd1619: dataIn2 = 32'd63; 
32'd1620: dataIn2 = 32'd89; 
32'd1621: dataIn2 = 32'd41; 
32'd1622: dataIn2 = 32'd52; 
32'd1623: dataIn2 = 32'd78; 
32'd1624: dataIn2 = 32'd100; 
32'd1625: dataIn2 = 32'd3; 
32'd1626: dataIn2 = 32'd75; 
32'd1627: dataIn2 = 32'd6; 
32'd1628: dataIn2 = 32'd79; 
32'd1629: dataIn2 = 32'd0; 
32'd1630: dataIn2 = 32'd18; 
32'd1631: dataIn2 = 32'd24; 
32'd1632: dataIn2 = 32'd42; 
32'd1633: dataIn2 = 32'd43; 
32'd1634: dataIn2 = 32'd3; 
32'd1635: dataIn2 = 32'd100; 
32'd1636: dataIn2 = 32'd28; 
32'd1637: dataIn2 = 32'd81; 
32'd1638: dataIn2 = 32'd21; 
32'd1639: dataIn2 = 32'd9; 
32'd1640: dataIn2 = 32'd54; 
32'd1641: dataIn2 = 32'd33; 
32'd1642: dataIn2 = 32'd97; 
32'd1643: dataIn2 = 32'd52; 
32'd1644: dataIn2 = 32'd24; 
32'd1645: dataIn2 = 32'd73; 
32'd1646: dataIn2 = 32'd12; 
32'd1647: dataIn2 = 32'd65; 
32'd1648: dataIn2 = 32'd23; 
32'd1649: dataIn2 = 32'd42; 
32'd1650: dataIn2 = 32'd59; 
32'd1651: dataIn2 = 32'd31; 
32'd1652: dataIn2 = 32'd84; 
32'd1653: dataIn2 = 32'd26; 
32'd1654: dataIn2 = 32'd27; 
32'd1655: dataIn2 = 32'd2; 
32'd1656: dataIn2 = 32'd77; 
32'd1657: dataIn2 = 32'd57; 
32'd1658: dataIn2 = 32'd1; 
32'd1659: dataIn2 = 32'd10; 
32'd1660: dataIn2 = 32'd28; 
32'd1661: dataIn2 = 32'd28; 
32'd1662: dataIn2 = 32'd61; 
32'd1663: dataIn2 = 32'd17; 
32'd1664: dataIn2 = 32'd78; 
32'd1665: dataIn2 = 32'd1; 
32'd1666: dataIn2 = 32'd40; 
32'd1667: dataIn2 = 32'd78; 
32'd1668: dataIn2 = 32'd52; 
32'd1669: dataIn2 = 32'd32; 
32'd1670: dataIn2 = 32'd92; 
32'd1671: dataIn2 = 32'd10; 
32'd1672: dataIn2 = 32'd67; 
32'd1673: dataIn2 = 32'd67; 
32'd1674: dataIn2 = 32'd11; 
32'd1675: dataIn2 = 32'd43; 
32'd1676: dataIn2 = 32'd51; 
32'd1677: dataIn2 = 32'd58; 
32'd1678: dataIn2 = 32'd80; 
32'd1679: dataIn2 = 32'd67; 
32'd1680: dataIn2 = 32'd37; 
32'd1681: dataIn2 = 32'd13; 
32'd1682: dataIn2 = 32'd94; 
32'd1683: dataIn2 = 32'd98; 
32'd1684: dataIn2 = 32'd74; 
32'd1685: dataIn2 = 32'd71; 
32'd1686: dataIn2 = 32'd95; 
32'd1687: dataIn2 = 32'd63; 
32'd1688: dataIn2 = 32'd59; 
32'd1689: dataIn2 = 32'd37; 
32'd1690: dataIn2 = 32'd95; 
32'd1691: dataIn2 = 32'd17; 
32'd1692: dataIn2 = 32'd2; 
32'd1693: dataIn2 = 32'd12; 
32'd1694: dataIn2 = 32'd39; 
32'd1695: dataIn2 = 32'd32; 
32'd1696: dataIn2 = 32'd87; 
32'd1697: dataIn2 = 32'd79; 
32'd1698: dataIn2 = 32'd75; 
32'd1699: dataIn2 = 32'd57; 
32'd1700: dataIn2 = 32'd14; 
32'd1701: dataIn2 = 32'd39; 
32'd1702: dataIn2 = 32'd82; 
32'd1703: dataIn2 = 32'd76; 
32'd1704: dataIn2 = 32'd77; 
32'd1705: dataIn2 = 32'd13; 
32'd1706: dataIn2 = 32'd75; 
32'd1707: dataIn2 = 32'd32; 
32'd1708: dataIn2 = 32'd89; 
32'd1709: dataIn2 = 32'd59; 
32'd1710: dataIn2 = 32'd55; 
32'd1711: dataIn2 = 32'd93; 
32'd1712: dataIn2 = 32'd21; 
32'd1713: dataIn2 = 32'd59; 
32'd1714: dataIn2 = 32'd56; 
32'd1715: dataIn2 = 32'd57; 
32'd1716: dataIn2 = 32'd28; 
32'd1717: dataIn2 = 32'd66; 
32'd1718: dataIn2 = 32'd52; 
32'd1719: dataIn2 = 32'd6; 
32'd1720: dataIn2 = 32'd97; 
32'd1721: dataIn2 = 32'd34; 
32'd1722: dataIn2 = 32'd71; 
32'd1723: dataIn2 = 32'd94; 
32'd1724: dataIn2 = 32'd88; 
32'd1725: dataIn2 = 32'd42; 
32'd1726: dataIn2 = 32'd73; 
32'd1727: dataIn2 = 32'd0; 
32'd1728: dataIn2 = 32'd76; 
32'd1729: dataIn2 = 32'd20; 
32'd1730: dataIn2 = 32'd76; 
32'd1731: dataIn2 = 32'd52; 
32'd1732: dataIn2 = 32'd34; 
32'd1733: dataIn2 = 32'd91; 
32'd1734: dataIn2 = 32'd77; 
32'd1735: dataIn2 = 32'd16; 
32'd1736: dataIn2 = 32'd88; 
32'd1737: dataIn2 = 32'd64; 
32'd1738: dataIn2 = 32'd23; 
32'd1739: dataIn2 = 32'd30; 
32'd1740: dataIn2 = 32'd99; 
32'd1741: dataIn2 = 32'd34; 
32'd1742: dataIn2 = 32'd0; 
32'd1743: dataIn2 = 32'd53; 
32'd1744: dataIn2 = 32'd51; 
32'd1745: dataIn2 = 32'd46; 
32'd1746: dataIn2 = 32'd78; 
32'd1747: dataIn2 = 32'd94; 
32'd1748: dataIn2 = 32'd58; 
32'd1749: dataIn2 = 32'd82; 
32'd1750: dataIn2 = 32'd30; 
32'd1751: dataIn2 = 32'd38; 
32'd1752: dataIn2 = 32'd87; 
32'd1753: dataIn2 = 32'd23; 
32'd1754: dataIn2 = 32'd17; 
32'd1755: dataIn2 = 32'd73; 
32'd1756: dataIn2 = 32'd21; 
32'd1757: dataIn2 = 32'd72; 
32'd1758: dataIn2 = 32'd57; 
32'd1759: dataIn2 = 32'd12; 
32'd1760: dataIn2 = 32'd97; 
32'd1761: dataIn2 = 32'd70; 
32'd1762: dataIn2 = 32'd19; 
32'd1763: dataIn2 = 32'd41; 
32'd1764: dataIn2 = 32'd65; 
32'd1765: dataIn2 = 32'd99; 
32'd1766: dataIn2 = 32'd45; 
32'd1767: dataIn2 = 32'd69; 
32'd1768: dataIn2 = 32'd39; 
32'd1769: dataIn2 = 32'd84; 
32'd1770: dataIn2 = 32'd43; 
32'd1771: dataIn2 = 32'd86; 
32'd1772: dataIn2 = 32'd4; 
32'd1773: dataIn2 = 32'd65; 
32'd1774: dataIn2 = 32'd43; 
32'd1775: dataIn2 = 32'd18; 
32'd1776: dataIn2 = 32'd20; 
32'd1777: dataIn2 = 32'd10; 
32'd1778: dataIn2 = 32'd15; 
32'd1779: dataIn2 = 32'd71; 
32'd1780: dataIn2 = 32'd16; 
32'd1781: dataIn2 = 32'd83; 
32'd1782: dataIn2 = 32'd23; 
32'd1783: dataIn2 = 32'd31; 
32'd1784: dataIn2 = 32'd43; 
32'd1785: dataIn2 = 32'd57; 
32'd1786: dataIn2 = 32'd22; 
32'd1787: dataIn2 = 32'd1; 
32'd1788: dataIn2 = 32'd16; 
32'd1789: dataIn2 = 32'd34; 
32'd1790: dataIn2 = 32'd87; 
32'd1791: dataIn2 = 32'd53; 
32'd1792: dataIn2 = 32'd52; 
32'd1793: dataIn2 = 32'd44; 
32'd1794: dataIn2 = 32'd33; 
32'd1795: dataIn2 = 32'd34; 
32'd1796: dataIn2 = 32'd18; 
32'd1797: dataIn2 = 32'd66; 
32'd1798: dataIn2 = 32'd28; 
32'd1799: dataIn2 = 32'd0; 
32'd1800: dataIn2 = 32'd65; 
32'd1801: dataIn2 = 32'd15; 
32'd1802: dataIn2 = 32'd3; 
32'd1803: dataIn2 = 32'd94; 
32'd1804: dataIn2 = 32'd24; 
32'd1805: dataIn2 = 32'd92; 
32'd1806: dataIn2 = 32'd9; 
32'd1807: dataIn2 = 32'd27; 
32'd1808: dataIn2 = 32'd1; 
32'd1809: dataIn2 = 32'd53; 
32'd1810: dataIn2 = 32'd64; 
32'd1811: dataIn2 = 32'd95; 
32'd1812: dataIn2 = 32'd67; 
32'd1813: dataIn2 = 32'd27; 
32'd1814: dataIn2 = 32'd9; 
32'd1815: dataIn2 = 32'd20; 
32'd1816: dataIn2 = 32'd29; 
32'd1817: dataIn2 = 32'd70; 
32'd1818: dataIn2 = 32'd1; 
32'd1819: dataIn2 = 32'd65; 
32'd1820: dataIn2 = 32'd34; 
32'd1821: dataIn2 = 32'd44; 
32'd1822: dataIn2 = 32'd100; 
32'd1823: dataIn2 = 32'd20; 
32'd1824: dataIn2 = 32'd11; 
32'd1825: dataIn2 = 32'd89; 
32'd1826: dataIn2 = 32'd62; 
32'd1827: dataIn2 = 32'd48; 
32'd1828: dataIn2 = 32'd81; 
32'd1829: dataIn2 = 32'd38; 
32'd1830: dataIn2 = 32'd75; 
32'd1831: dataIn2 = 32'd33; 
32'd1832: dataIn2 = 32'd57; 
32'd1833: dataIn2 = 32'd89; 
32'd1834: dataIn2 = 32'd1; 
32'd1835: dataIn2 = 32'd32; 
32'd1836: dataIn2 = 32'd8; 
32'd1837: dataIn2 = 32'd56; 
32'd1838: dataIn2 = 32'd100; 
32'd1839: dataIn2 = 32'd53; 
32'd1840: dataIn2 = 32'd14; 
32'd1841: dataIn2 = 32'd56; 
32'd1842: dataIn2 = 32'd40; 
32'd1843: dataIn2 = 32'd12; 
32'd1844: dataIn2 = 32'd33; 
32'd1845: dataIn2 = 32'd6; 
32'd1846: dataIn2 = 32'd69; 
32'd1847: dataIn2 = 32'd1; 
32'd1848: dataIn2 = 32'd48; 
32'd1849: dataIn2 = 32'd70; 
32'd1850: dataIn2 = 32'd95; 
32'd1851: dataIn2 = 32'd46; 
32'd1852: dataIn2 = 32'd22; 
32'd1853: dataIn2 = 32'd49; 
32'd1854: dataIn2 = 32'd91; 
32'd1855: dataIn2 = 32'd14; 
32'd1856: dataIn2 = 32'd56; 
32'd1857: dataIn2 = 32'd60; 
32'd1858: dataIn2 = 32'd93; 
32'd1859: dataIn2 = 32'd72; 
32'd1860: dataIn2 = 32'd67; 
32'd1861: dataIn2 = 32'd55; 
32'd1862: dataIn2 = 32'd6; 
32'd1863: dataIn2 = 32'd35; 
32'd1864: dataIn2 = 32'd86; 
32'd1865: dataIn2 = 32'd34; 
32'd1866: dataIn2 = 32'd24; 
32'd1867: dataIn2 = 32'd22; 
32'd1868: dataIn2 = 32'd47; 
32'd1869: dataIn2 = 32'd90; 
32'd1870: dataIn2 = 32'd5; 
32'd1871: dataIn2 = 32'd14; 
32'd1872: dataIn2 = 32'd61; 
32'd1873: dataIn2 = 32'd21; 
32'd1874: dataIn2 = 32'd56; 
32'd1875: dataIn2 = 32'd64; 
32'd1876: dataIn2 = 32'd82; 
32'd1877: dataIn2 = 32'd64; 
32'd1878: dataIn2 = 32'd28; 
32'd1879: dataIn2 = 32'd27; 
32'd1880: dataIn2 = 32'd97; 
32'd1881: dataIn2 = 32'd61; 
32'd1882: dataIn2 = 32'd54; 
32'd1883: dataIn2 = 32'd77; 
32'd1884: dataIn2 = 32'd2; 
32'd1885: dataIn2 = 32'd34; 
32'd1886: dataIn2 = 32'd66; 
32'd1887: dataIn2 = 32'd80; 
32'd1888: dataIn2 = 32'd11; 
32'd1889: dataIn2 = 32'd68; 
32'd1890: dataIn2 = 32'd50; 
32'd1891: dataIn2 = 32'd32; 
32'd1892: dataIn2 = 32'd53; 
32'd1893: dataIn2 = 32'd75; 
32'd1894: dataIn2 = 32'd29; 
32'd1895: dataIn2 = 32'd98; 
32'd1896: dataIn2 = 32'd33; 
32'd1897: dataIn2 = 32'd37; 
32'd1898: dataIn2 = 32'd45; 
32'd1899: dataIn2 = 32'd30; 
32'd1900: dataIn2 = 32'd2; 
32'd1901: dataIn2 = 32'd27; 
32'd1902: dataIn2 = 32'd93; 
32'd1903: dataIn2 = 32'd65; 
32'd1904: dataIn2 = 32'd28; 
32'd1905: dataIn2 = 32'd11; 
32'd1906: dataIn2 = 32'd25; 
32'd1907: dataIn2 = 32'd67; 
32'd1908: dataIn2 = 32'd96; 
32'd1909: dataIn2 = 32'd80; 
32'd1910: dataIn2 = 32'd98; 
32'd1911: dataIn2 = 32'd9; 
32'd1912: dataIn2 = 32'd8; 
32'd1913: dataIn2 = 32'd41; 
32'd1914: dataIn2 = 32'd100; 
32'd1915: dataIn2 = 32'd65; 
32'd1916: dataIn2 = 32'd19; 
32'd1917: dataIn2 = 32'd21; 
32'd1918: dataIn2 = 32'd84; 
32'd1919: dataIn2 = 32'd86; 
32'd1920: dataIn2 = 32'd61; 
32'd1921: dataIn2 = 32'd87; 
32'd1922: dataIn2 = 32'd10; 
32'd1923: dataIn2 = 32'd29; 
32'd1924: dataIn2 = 32'd92; 
32'd1925: dataIn2 = 32'd16; 
32'd1926: dataIn2 = 32'd18; 
32'd1927: dataIn2 = 32'd87; 
32'd1928: dataIn2 = 32'd48; 
32'd1929: dataIn2 = 32'd25; 
32'd1930: dataIn2 = 32'd92; 
32'd1931: dataIn2 = 32'd3; 
32'd1932: dataIn2 = 32'd98; 
32'd1933: dataIn2 = 32'd33; 
32'd1934: dataIn2 = 32'd16; 
32'd1935: dataIn2 = 32'd20; 
32'd1936: dataIn2 = 32'd1; 
32'd1937: dataIn2 = 32'd93; 
32'd1938: dataIn2 = 32'd12; 
32'd1939: dataIn2 = 32'd20; 
32'd1940: dataIn2 = 32'd30; 
32'd1941: dataIn2 = 32'd76; 
32'd1942: dataIn2 = 32'd29; 
32'd1943: dataIn2 = 32'd98; 
32'd1944: dataIn2 = 32'd69; 
32'd1945: dataIn2 = 32'd59; 
32'd1946: dataIn2 = 32'd29; 
32'd1947: dataIn2 = 32'd53; 
32'd1948: dataIn2 = 32'd32; 
32'd1949: dataIn2 = 32'd88; 
32'd1950: dataIn2 = 32'd6; 
32'd1951: dataIn2 = 32'd54; 
32'd1952: dataIn2 = 32'd66; 
32'd1953: dataIn2 = 32'd89; 
32'd1954: dataIn2 = 32'd25; 
32'd1955: dataIn2 = 32'd75; 
32'd1956: dataIn2 = 32'd100; 
32'd1957: dataIn2 = 32'd22; 
32'd1958: dataIn2 = 32'd24; 
32'd1959: dataIn2 = 32'd47; 
32'd1960: dataIn2 = 32'd55; 
32'd1961: dataIn2 = 32'd56; 
32'd1962: dataIn2 = 32'd6; 
32'd1963: dataIn2 = 32'd88; 
32'd1964: dataIn2 = 32'd10; 
32'd1965: dataIn2 = 32'd53; 
32'd1966: dataIn2 = 32'd87; 
32'd1967: dataIn2 = 32'd29; 
32'd1968: dataIn2 = 32'd53; 
32'd1969: dataIn2 = 32'd16; 
32'd1970: dataIn2 = 32'd74; 
32'd1971: dataIn2 = 32'd87; 
32'd1972: dataIn2 = 32'd4; 
32'd1973: dataIn2 = 32'd64; 
32'd1974: dataIn2 = 32'd77; 
32'd1975: dataIn2 = 32'd33; 
32'd1976: dataIn2 = 32'd90; 
32'd1977: dataIn2 = 32'd38; 
32'd1978: dataIn2 = 32'd31; 
32'd1979: dataIn2 = 32'd27; 
32'd1980: dataIn2 = 32'd53; 
32'd1981: dataIn2 = 32'd83; 
32'd1982: dataIn2 = 32'd95; 
32'd1983: dataIn2 = 32'd96; 
32'd1984: dataIn2 = 32'd63; 
32'd1985: dataIn2 = 32'd72; 
32'd1986: dataIn2 = 32'd86; 
32'd1987: dataIn2 = 32'd5; 
32'd1988: dataIn2 = 32'd29; 
32'd1989: dataIn2 = 32'd64; 
32'd1990: dataIn2 = 32'd0; 
32'd1991: dataIn2 = 32'd49; 
32'd1992: dataIn2 = 32'd91; 
32'd1993: dataIn2 = 32'd83; 
32'd1994: dataIn2 = 32'd6; 
32'd1995: dataIn2 = 32'd27; 
32'd1996: dataIn2 = 32'd77; 
32'd1997: dataIn2 = 32'd68; 
32'd1998: dataIn2 = 32'd92; 
32'd1999: dataIn2 = 32'd54; 
32'd2000: dataIn2 = 32'd43; 
32'd2001: dataIn2 = 32'd92; 
32'd2002: dataIn2 = 32'd30; 
32'd2003: dataIn2 = 32'd82; 
32'd2004: dataIn2 = 32'd42; 
32'd2005: dataIn2 = 32'd97; 
32'd2006: dataIn2 = 32'd87; 
32'd2007: dataIn2 = 32'd14; 
32'd2008: dataIn2 = 32'd12; 
32'd2009: dataIn2 = 32'd63; 
32'd2010: dataIn2 = 32'd29; 
32'd2011: dataIn2 = 32'd57; 
32'd2012: dataIn2 = 32'd64; 
32'd2013: dataIn2 = 32'd74; 
32'd2014: dataIn2 = 32'd100; 
32'd2015: dataIn2 = 32'd68; 
32'd2016: dataIn2 = 32'd96; 
32'd2017: dataIn2 = 32'd57; 
32'd2018: dataIn2 = 32'd47; 
32'd2019: dataIn2 = 32'd52; 
32'd2020: dataIn2 = 32'd30; 
32'd2021: dataIn2 = 32'd30; 
32'd2022: dataIn2 = 32'd87; 
32'd2023: dataIn2 = 32'd30; 
32'd2024: dataIn2 = 32'd9; 
32'd2025: dataIn2 = 32'd81; 
32'd2026: dataIn2 = 32'd98; 
32'd2027: dataIn2 = 32'd38; 
32'd2028: dataIn2 = 32'd51; 
32'd2029: dataIn2 = 32'd81; 
32'd2030: dataIn2 = 32'd49; 
32'd2031: dataIn2 = 32'd48; 
32'd2032: dataIn2 = 32'd25; 
32'd2033: dataIn2 = 32'd61; 
32'd2034: dataIn2 = 32'd68; 
32'd2035: dataIn2 = 32'd23; 
32'd2036: dataIn2 = 32'd87; 
32'd2037: dataIn2 = 32'd13; 
32'd2038: dataIn2 = 32'd31; 
32'd2039: dataIn2 = 32'd48; 
32'd2040: dataIn2 = 32'd4; 
32'd2041: dataIn2 = 32'd43; 
32'd2042: dataIn2 = 32'd38; 
32'd2043: dataIn2 = 32'd87; 
32'd2044: dataIn2 = 32'd28; 
32'd2045: dataIn2 = 32'd45; 
32'd2046: dataIn2 = 32'd34; 
32'd2047: dataIn2 = 32'd15; 
32'd2048: dataIn2 = 32'd46; 
32'd2049: dataIn2 = 32'd55; 
32'd2050: dataIn2 = 32'd43; 
32'd2051: dataIn2 = 32'd95; 
32'd2052: dataIn2 = 32'd2; 
32'd2053: dataIn2 = 32'd27; 
32'd2054: dataIn2 = 32'd21; 
32'd2055: dataIn2 = 32'd86; 
32'd2056: dataIn2 = 32'd89; 
32'd2057: dataIn2 = 32'd86; 
32'd2058: dataIn2 = 32'd73; 
32'd2059: dataIn2 = 32'd89; 
32'd2060: dataIn2 = 32'd24; 
32'd2061: dataIn2 = 32'd40; 
32'd2062: dataIn2 = 32'd99; 
32'd2063: dataIn2 = 32'd62; 
32'd2064: dataIn2 = 32'd33; 
32'd2065: dataIn2 = 32'd3; 
32'd2066: dataIn2 = 32'd41; 
32'd2067: dataIn2 = 32'd22; 
32'd2068: dataIn2 = 32'd1; 
32'd2069: dataIn2 = 32'd40; 
32'd2070: dataIn2 = 32'd18; 
32'd2071: dataIn2 = 32'd8; 
32'd2072: dataIn2 = 32'd83; 
32'd2073: dataIn2 = 32'd18; 
32'd2074: dataIn2 = 32'd86; 
32'd2075: dataIn2 = 32'd98; 
32'd2076: dataIn2 = 32'd82; 
32'd2077: dataIn2 = 32'd56; 
32'd2078: dataIn2 = 32'd0; 
32'd2079: dataIn2 = 32'd48; 
32'd2080: dataIn2 = 32'd57; 
32'd2081: dataIn2 = 32'd3; 
32'd2082: dataIn2 = 32'd74; 
32'd2083: dataIn2 = 32'd94; 
32'd2084: dataIn2 = 32'd23; 
32'd2085: dataIn2 = 32'd20; 
32'd2086: dataIn2 = 32'd24; 
32'd2087: dataIn2 = 32'd1; 
32'd2088: dataIn2 = 32'd84; 
32'd2089: dataIn2 = 32'd3; 
32'd2090: dataIn2 = 32'd91; 
32'd2091: dataIn2 = 32'd1; 
32'd2092: dataIn2 = 32'd61; 
32'd2093: dataIn2 = 32'd72; 
32'd2094: dataIn2 = 32'd50; 
32'd2095: dataIn2 = 32'd83; 
32'd2096: dataIn2 = 32'd27; 
32'd2097: dataIn2 = 32'd92; 
32'd2098: dataIn2 = 32'd46; 
32'd2099: dataIn2 = 32'd2; 
32'd2100: dataIn2 = 32'd33; 
32'd2101: dataIn2 = 32'd19; 
32'd2102: dataIn2 = 32'd79; 
32'd2103: dataIn2 = 32'd27; 
32'd2104: dataIn2 = 32'd28; 
32'd2105: dataIn2 = 32'd31; 
32'd2106: dataIn2 = 32'd14; 
32'd2107: dataIn2 = 32'd32; 
32'd2108: dataIn2 = 32'd86; 
32'd2109: dataIn2 = 32'd32; 
32'd2110: dataIn2 = 32'd40; 
32'd2111: dataIn2 = 32'd88; 
32'd2112: dataIn2 = 32'd97; 
32'd2113: dataIn2 = 32'd0; 
32'd2114: dataIn2 = 32'd25; 
32'd2115: dataIn2 = 32'd50; 
32'd2116: dataIn2 = 32'd63; 
32'd2117: dataIn2 = 32'd70; 
32'd2118: dataIn2 = 32'd18; 
32'd2119: dataIn2 = 32'd16; 
32'd2120: dataIn2 = 32'd80; 
32'd2121: dataIn2 = 32'd14; 
32'd2122: dataIn2 = 32'd89; 
32'd2123: dataIn2 = 32'd45; 
32'd2124: dataIn2 = 32'd55; 
32'd2125: dataIn2 = 32'd86; 
32'd2126: dataIn2 = 32'd54; 
32'd2127: dataIn2 = 32'd20; 
32'd2128: dataIn2 = 32'd18; 
32'd2129: dataIn2 = 32'd68; 
32'd2130: dataIn2 = 32'd47; 
32'd2131: dataIn2 = 32'd29; 
32'd2132: dataIn2 = 32'd67; 
32'd2133: dataIn2 = 32'd56; 
32'd2134: dataIn2 = 32'd39; 
32'd2135: dataIn2 = 32'd13; 
32'd2136: dataIn2 = 32'd37; 
32'd2137: dataIn2 = 32'd19; 
32'd2138: dataIn2 = 32'd64; 
32'd2139: dataIn2 = 32'd48; 
32'd2140: dataIn2 = 32'd73; 
32'd2141: dataIn2 = 32'd82; 
32'd2142: dataIn2 = 32'd17; 
32'd2143: dataIn2 = 32'd64; 
32'd2144: dataIn2 = 32'd94; 
32'd2145: dataIn2 = 32'd19; 
32'd2146: dataIn2 = 32'd45; 
32'd2147: dataIn2 = 32'd81; 
32'd2148: dataIn2 = 32'd29; 
32'd2149: dataIn2 = 32'd3; 
32'd2150: dataIn2 = 32'd7; 
32'd2151: dataIn2 = 32'd84; 
32'd2152: dataIn2 = 32'd93; 
32'd2153: dataIn2 = 32'd71; 
32'd2154: dataIn2 = 32'd23; 
32'd2155: dataIn2 = 32'd69; 
32'd2156: dataIn2 = 32'd30; 
32'd2157: dataIn2 = 32'd48; 
32'd2158: dataIn2 = 32'd55; 
32'd2159: dataIn2 = 32'd98; 
32'd2160: dataIn2 = 32'd33; 
32'd2161: dataIn2 = 32'd6; 
32'd2162: dataIn2 = 32'd16; 
32'd2163: dataIn2 = 32'd66; 
32'd2164: dataIn2 = 32'd29; 
32'd2165: dataIn2 = 32'd5; 
32'd2166: dataIn2 = 32'd68; 
32'd2167: dataIn2 = 32'd95; 
32'd2168: dataIn2 = 32'd71; 
32'd2169: dataIn2 = 32'd95; 
32'd2170: dataIn2 = 32'd91; 
32'd2171: dataIn2 = 32'd0; 
32'd2172: dataIn2 = 32'd2; 
32'd2173: dataIn2 = 32'd20; 
32'd2174: dataIn2 = 32'd52; 
32'd2175: dataIn2 = 32'd44; 
32'd2176: dataIn2 = 32'd9; 
32'd2177: dataIn2 = 32'd91; 
32'd2178: dataIn2 = 32'd67; 
32'd2179: dataIn2 = 32'd63; 
32'd2180: dataIn2 = 32'd5; 
32'd2181: dataIn2 = 32'd33; 
32'd2182: dataIn2 = 32'd29; 
32'd2183: dataIn2 = 32'd9; 
32'd2184: dataIn2 = 32'd22; 
32'd2185: dataIn2 = 32'd38; 
32'd2186: dataIn2 = 32'd5; 
32'd2187: dataIn2 = 32'd59; 
32'd2188: dataIn2 = 32'd96; 
32'd2189: dataIn2 = 32'd90; 
32'd2190: dataIn2 = 32'd92; 
32'd2191: dataIn2 = 32'd31; 
32'd2192: dataIn2 = 32'd16; 
32'd2193: dataIn2 = 32'd81; 
32'd2194: dataIn2 = 32'd12; 
32'd2195: dataIn2 = 32'd34; 
32'd2196: dataIn2 = 32'd96; 
32'd2197: dataIn2 = 32'd79; 
32'd2198: dataIn2 = 32'd70; 
32'd2199: dataIn2 = 32'd50; 
32'd2200: dataIn2 = 32'd7; 
32'd2201: dataIn2 = 32'd99; 
32'd2202: dataIn2 = 32'd63; 
32'd2203: dataIn2 = 32'd99; 
32'd2204: dataIn2 = 32'd33; 
32'd2205: dataIn2 = 32'd17; 
32'd2206: dataIn2 = 32'd86; 
32'd2207: dataIn2 = 32'd10; 
32'd2208: dataIn2 = 32'd66; 
32'd2209: dataIn2 = 32'd15; 
32'd2210: dataIn2 = 32'd85; 
32'd2211: dataIn2 = 32'd77; 
32'd2212: dataIn2 = 32'd71; 
32'd2213: dataIn2 = 32'd72; 
32'd2214: dataIn2 = 32'd40; 
32'd2215: dataIn2 = 32'd92; 
32'd2216: dataIn2 = 32'd78; 
32'd2217: dataIn2 = 32'd45; 
32'd2218: dataIn2 = 32'd35; 
32'd2219: dataIn2 = 32'd79; 
32'd2220: dataIn2 = 32'd28; 
32'd2221: dataIn2 = 32'd9; 
32'd2222: dataIn2 = 32'd78; 
32'd2223: dataIn2 = 32'd23; 
32'd2224: dataIn2 = 32'd88; 
32'd2225: dataIn2 = 32'd96; 
32'd2226: dataIn2 = 32'd12; 
32'd2227: dataIn2 = 32'd46; 
32'd2228: dataIn2 = 32'd41; 
32'd2229: dataIn2 = 32'd81; 
32'd2230: dataIn2 = 32'd60; 
32'd2231: dataIn2 = 32'd4; 
32'd2232: dataIn2 = 32'd4; 
32'd2233: dataIn2 = 32'd3; 
32'd2234: dataIn2 = 32'd26; 
32'd2235: dataIn2 = 32'd49; 
32'd2236: dataIn2 = 32'd23; 
32'd2237: dataIn2 = 32'd38; 
32'd2238: dataIn2 = 32'd62; 
32'd2239: dataIn2 = 32'd9; 
32'd2240: dataIn2 = 32'd73; 
32'd2241: dataIn2 = 32'd43; 
32'd2242: dataIn2 = 32'd45; 
32'd2243: dataIn2 = 32'd1; 
32'd2244: dataIn2 = 32'd41; 
32'd2245: dataIn2 = 32'd63; 
32'd2246: dataIn2 = 32'd79; 
32'd2247: dataIn2 = 32'd41; 
32'd2248: dataIn2 = 32'd75; 
32'd2249: dataIn2 = 32'd31; 
32'd2250: dataIn2 = 32'd26; 
32'd2251: dataIn2 = 32'd76; 
32'd2252: dataIn2 = 32'd0; 
32'd2253: dataIn2 = 32'd82; 
32'd2254: dataIn2 = 32'd1; 
32'd2255: dataIn2 = 32'd38; 
32'd2256: dataIn2 = 32'd17; 
32'd2257: dataIn2 = 32'd27; 
32'd2258: dataIn2 = 32'd10; 
32'd2259: dataIn2 = 32'd81; 
32'd2260: dataIn2 = 32'd62; 
32'd2261: dataIn2 = 32'd43; 
32'd2262: dataIn2 = 32'd17; 
32'd2263: dataIn2 = 32'd90; 
32'd2264: dataIn2 = 32'd26; 
32'd2265: dataIn2 = 32'd9; 
32'd2266: dataIn2 = 32'd40; 
32'd2267: dataIn2 = 32'd40; 
32'd2268: dataIn2 = 32'd34; 
32'd2269: dataIn2 = 32'd37; 
32'd2270: dataIn2 = 32'd49; 
32'd2271: dataIn2 = 32'd13; 
32'd2272: dataIn2 = 32'd23; 
32'd2273: dataIn2 = 32'd62; 
32'd2274: dataIn2 = 32'd70; 
32'd2275: dataIn2 = 32'd10; 
32'd2276: dataIn2 = 32'd3; 
32'd2277: dataIn2 = 32'd23; 
32'd2278: dataIn2 = 32'd75; 
32'd2279: dataIn2 = 32'd27; 
32'd2280: dataIn2 = 32'd84; 
32'd2281: dataIn2 = 32'd70; 
32'd2282: dataIn2 = 32'd88; 
32'd2283: dataIn2 = 32'd23; 
32'd2284: dataIn2 = 32'd96; 
32'd2285: dataIn2 = 32'd45; 
32'd2286: dataIn2 = 32'd91; 
32'd2287: dataIn2 = 32'd31; 
32'd2288: dataIn2 = 32'd60; 
32'd2289: dataIn2 = 32'd27; 
32'd2290: dataIn2 = 32'd77; 
32'd2291: dataIn2 = 32'd18; 
32'd2292: dataIn2 = 32'd80; 
32'd2293: dataIn2 = 32'd8; 
32'd2294: dataIn2 = 32'd21; 
32'd2295: dataIn2 = 32'd17; 
32'd2296: dataIn2 = 32'd18; 
32'd2297: dataIn2 = 32'd12; 
32'd2298: dataIn2 = 32'd13; 
32'd2299: dataIn2 = 32'd63; 
32'd2300: dataIn2 = 32'd13; 
32'd2301: dataIn2 = 32'd27; 
32'd2302: dataIn2 = 32'd15; 
32'd2303: dataIn2 = 32'd96; 
32'd2304: dataIn2 = 32'd53; 
32'd2305: dataIn2 = 32'd84; 
32'd2306: dataIn2 = 32'd31; 
32'd2307: dataIn2 = 32'd46; 
32'd2308: dataIn2 = 32'd53; 
32'd2309: dataIn2 = 32'd61; 
32'd2310: dataIn2 = 32'd49; 
32'd2311: dataIn2 = 32'd38; 
32'd2312: dataIn2 = 32'd32; 
32'd2313: dataIn2 = 32'd12; 
32'd2314: dataIn2 = 32'd71; 
32'd2315: dataIn2 = 32'd4; 
32'd2316: dataIn2 = 32'd18; 
32'd2317: dataIn2 = 32'd98; 
32'd2318: dataIn2 = 32'd27; 
32'd2319: dataIn2 = 32'd18; 
32'd2320: dataIn2 = 32'd79; 
32'd2321: dataIn2 = 32'd38; 
32'd2322: dataIn2 = 32'd59; 
32'd2323: dataIn2 = 32'd37; 
32'd2324: dataIn2 = 32'd59; 
32'd2325: dataIn2 = 32'd17; 
32'd2326: dataIn2 = 32'd58; 
32'd2327: dataIn2 = 32'd76; 
32'd2328: dataIn2 = 32'd10; 
32'd2329: dataIn2 = 32'd63; 
32'd2330: dataIn2 = 32'd65; 
32'd2331: dataIn2 = 32'd78; 
32'd2332: dataIn2 = 32'd73; 
32'd2333: dataIn2 = 32'd98; 
32'd2334: dataIn2 = 32'd68; 
32'd2335: dataIn2 = 32'd53; 
32'd2336: dataIn2 = 32'd27; 
32'd2337: dataIn2 = 32'd92; 
32'd2338: dataIn2 = 32'd38; 
32'd2339: dataIn2 = 32'd73; 
32'd2340: dataIn2 = 32'd59; 
32'd2341: dataIn2 = 32'd75; 
32'd2342: dataIn2 = 32'd42; 
32'd2343: dataIn2 = 32'd13; 
32'd2344: dataIn2 = 32'd25; 
32'd2345: dataIn2 = 32'd75; 
32'd2346: dataIn2 = 32'd16; 
32'd2347: dataIn2 = 32'd85; 
32'd2348: dataIn2 = 32'd23; 
32'd2349: dataIn2 = 32'd99; 
32'd2350: dataIn2 = 32'd87; 
32'd2351: dataIn2 = 32'd40; 
32'd2352: dataIn2 = 32'd26; 
32'd2353: dataIn2 = 32'd7; 
32'd2354: dataIn2 = 32'd14; 
32'd2355: dataIn2 = 32'd80; 
32'd2356: dataIn2 = 32'd37; 
32'd2357: dataIn2 = 32'd59; 
32'd2358: dataIn2 = 32'd38; 
32'd2359: dataIn2 = 32'd51; 
32'd2360: dataIn2 = 32'd78; 
32'd2361: dataIn2 = 32'd11; 
32'd2362: dataIn2 = 32'd93; 
32'd2363: dataIn2 = 32'd14; 
32'd2364: dataIn2 = 32'd84; 
32'd2365: dataIn2 = 32'd84; 
32'd2366: dataIn2 = 32'd55; 
32'd2367: dataIn2 = 32'd70; 
32'd2368: dataIn2 = 32'd63; 
32'd2369: dataIn2 = 32'd98; 
32'd2370: dataIn2 = 32'd52; 
32'd2371: dataIn2 = 32'd22; 
32'd2372: dataIn2 = 32'd1; 
32'd2373: dataIn2 = 32'd56; 
32'd2374: dataIn2 = 32'd59; 
32'd2375: dataIn2 = 32'd89; 
32'd2376: dataIn2 = 32'd28; 
32'd2377: dataIn2 = 32'd15; 
32'd2378: dataIn2 = 32'd76; 
32'd2379: dataIn2 = 32'd80; 
32'd2380: dataIn2 = 32'd49; 
32'd2381: dataIn2 = 32'd88; 
32'd2382: dataIn2 = 32'd3; 
32'd2383: dataIn2 = 32'd52; 
32'd2384: dataIn2 = 32'd45; 
32'd2385: dataIn2 = 32'd70; 
32'd2386: dataIn2 = 32'd81; 
32'd2387: dataIn2 = 32'd58; 
32'd2388: dataIn2 = 32'd23; 
32'd2389: dataIn2 = 32'd54; 
32'd2390: dataIn2 = 32'd42; 
32'd2391: dataIn2 = 32'd1; 
32'd2392: dataIn2 = 32'd94; 
32'd2393: dataIn2 = 32'd29; 
32'd2394: dataIn2 = 32'd16; 
32'd2395: dataIn2 = 32'd19; 
32'd2396: dataIn2 = 32'd40; 
32'd2397: dataIn2 = 32'd1; 
32'd2398: dataIn2 = 32'd89; 
32'd2399: dataIn2 = 32'd69; 
32'd2400: dataIn2 = 32'd75; 
32'd2401: dataIn2 = 32'd81; 
32'd2402: dataIn2 = 32'd72; 
32'd2403: dataIn2 = 32'd56; 
32'd2404: dataIn2 = 32'd43; 
32'd2405: dataIn2 = 32'd79; 
32'd2406: dataIn2 = 32'd73; 
32'd2407: dataIn2 = 32'd59; 
32'd2408: dataIn2 = 32'd60; 
32'd2409: dataIn2 = 32'd43; 
32'd2410: dataIn2 = 32'd96; 
32'd2411: dataIn2 = 32'd22; 
32'd2412: dataIn2 = 32'd27; 
32'd2413: dataIn2 = 32'd88; 
32'd2414: dataIn2 = 32'd14; 
32'd2415: dataIn2 = 32'd84; 
32'd2416: dataIn2 = 32'd67; 
32'd2417: dataIn2 = 32'd74; 
32'd2418: dataIn2 = 32'd20; 
32'd2419: dataIn2 = 32'd2; 
32'd2420: dataIn2 = 32'd82; 
32'd2421: dataIn2 = 32'd93; 
32'd2422: dataIn2 = 32'd55; 
32'd2423: dataIn2 = 32'd30; 
32'd2424: dataIn2 = 32'd55; 
32'd2425: dataIn2 = 32'd82; 
32'd2426: dataIn2 = 32'd56; 
32'd2427: dataIn2 = 32'd30; 
32'd2428: dataIn2 = 32'd27; 
32'd2429: dataIn2 = 32'd50; 
32'd2430: dataIn2 = 32'd34; 
32'd2431: dataIn2 = 32'd24; 
32'd2432: dataIn2 = 32'd9; 
32'd2433: dataIn2 = 32'd21; 
32'd2434: dataIn2 = 32'd5; 
32'd2435: dataIn2 = 32'd95; 
32'd2436: dataIn2 = 32'd83; 
32'd2437: dataIn2 = 32'd72; 
32'd2438: dataIn2 = 32'd50; 
32'd2439: dataIn2 = 32'd72; 
32'd2440: dataIn2 = 32'd6; 
32'd2441: dataIn2 = 32'd39; 
32'd2442: dataIn2 = 32'd89; 
32'd2443: dataIn2 = 32'd37; 
32'd2444: dataIn2 = 32'd36; 
32'd2445: dataIn2 = 32'd91; 
32'd2446: dataIn2 = 32'd16; 
32'd2447: dataIn2 = 32'd27; 
32'd2448: dataIn2 = 32'd82; 
32'd2449: dataIn2 = 32'd13; 
32'd2450: dataIn2 = 32'd18; 
32'd2451: dataIn2 = 32'd40; 
32'd2452: dataIn2 = 32'd74; 
32'd2453: dataIn2 = 32'd52; 
32'd2454: dataIn2 = 32'd27; 
32'd2455: dataIn2 = 32'd33; 
32'd2456: dataIn2 = 32'd79; 
32'd2457: dataIn2 = 32'd90; 
32'd2458: dataIn2 = 32'd19; 
32'd2459: dataIn2 = 32'd49; 
32'd2460: dataIn2 = 32'd57; 
32'd2461: dataIn2 = 32'd34; 
32'd2462: dataIn2 = 32'd25; 
32'd2463: dataIn2 = 32'd95; 
32'd2464: dataIn2 = 32'd65; 
32'd2465: dataIn2 = 32'd66; 
32'd2466: dataIn2 = 32'd53; 
32'd2467: dataIn2 = 32'd6; 
32'd2468: dataIn2 = 32'd57; 
32'd2469: dataIn2 = 32'd31; 
32'd2470: dataIn2 = 32'd12; 
32'd2471: dataIn2 = 32'd7; 
32'd2472: dataIn2 = 32'd42; 
32'd2473: dataIn2 = 32'd0; 
32'd2474: dataIn2 = 32'd72; 
32'd2475: dataIn2 = 32'd13; 
32'd2476: dataIn2 = 32'd45; 
32'd2477: dataIn2 = 32'd59; 
32'd2478: dataIn2 = 32'd0; 
32'd2479: dataIn2 = 32'd15; 
32'd2480: dataIn2 = 32'd51; 
32'd2481: dataIn2 = 32'd41; 
32'd2482: dataIn2 = 32'd51; 
32'd2483: dataIn2 = 32'd91; 
32'd2484: dataIn2 = 32'd2; 
32'd2485: dataIn2 = 32'd35; 
32'd2486: dataIn2 = 32'd98; 
32'd2487: dataIn2 = 32'd7; 
32'd2488: dataIn2 = 32'd85; 
32'd2489: dataIn2 = 32'd46; 
32'd2490: dataIn2 = 32'd94; 
32'd2491: dataIn2 = 32'd12; 
32'd2492: dataIn2 = 32'd62; 
32'd2493: dataIn2 = 32'd34; 
32'd2494: dataIn2 = 32'd88; 
32'd2495: dataIn2 = 32'd6; 
32'd2496: dataIn2 = 32'd87; 
32'd2497: dataIn2 = 32'd33; 
32'd2498: dataIn2 = 32'd84; 
32'd2499: dataIn2 = 32'd47; 
32'd2500: dataIn2 = 32'd41; 
32'd2501: dataIn2 = 32'd9; 
32'd2502: dataIn2 = 32'd56; 
32'd2503: dataIn2 = 32'd42; 
32'd2504: dataIn2 = 32'd80; 
32'd2505: dataIn2 = 32'd82; 
32'd2506: dataIn2 = 32'd98; 
32'd2507: dataIn2 = 32'd38; 
32'd2508: dataIn2 = 32'd40; 
32'd2509: dataIn2 = 32'd85; 
32'd2510: dataIn2 = 32'd7; 
32'd2511: dataIn2 = 32'd8; 
32'd2512: dataIn2 = 32'd36; 
32'd2513: dataIn2 = 32'd90; 
32'd2514: dataIn2 = 32'd43; 
32'd2515: dataIn2 = 32'd8; 
32'd2516: dataIn2 = 32'd17; 
32'd2517: dataIn2 = 32'd13; 
32'd2518: dataIn2 = 32'd43; 
32'd2519: dataIn2 = 32'd27; 
32'd2520: dataIn2 = 32'd79; 
32'd2521: dataIn2 = 32'd80; 
32'd2522: dataIn2 = 32'd9; 
32'd2523: dataIn2 = 32'd93; 
32'd2524: dataIn2 = 32'd42; 
32'd2525: dataIn2 = 32'd49; 
32'd2526: dataIn2 = 32'd81; 
32'd2527: dataIn2 = 32'd37; 
32'd2528: dataIn2 = 32'd39; 
32'd2529: dataIn2 = 32'd25; 
32'd2530: dataIn2 = 32'd89; 
32'd2531: dataIn2 = 32'd29; 
32'd2532: dataIn2 = 32'd41; 
32'd2533: dataIn2 = 32'd53; 
32'd2534: dataIn2 = 32'd92; 
32'd2535: dataIn2 = 32'd14; 
32'd2536: dataIn2 = 32'd48; 
32'd2537: dataIn2 = 32'd84; 
32'd2538: dataIn2 = 32'd57; 
32'd2539: dataIn2 = 32'd66; 
32'd2540: dataIn2 = 32'd72; 
32'd2541: dataIn2 = 32'd86; 
32'd2542: dataIn2 = 32'd39; 
32'd2543: dataIn2 = 32'd62; 
32'd2544: dataIn2 = 32'd92; 
32'd2545: dataIn2 = 32'd81; 
32'd2546: dataIn2 = 32'd68; 
32'd2547: dataIn2 = 32'd32; 
32'd2548: dataIn2 = 32'd68; 
32'd2549: dataIn2 = 32'd21; 
32'd2550: dataIn2 = 32'd38; 
32'd2551: dataIn2 = 32'd49; 
32'd2552: dataIn2 = 32'd67; 
32'd2553: dataIn2 = 32'd9; 
32'd2554: dataIn2 = 32'd94; 
32'd2555: dataIn2 = 32'd66; 
32'd2556: dataIn2 = 32'd70; 
32'd2557: dataIn2 = 32'd12; 
32'd2558: dataIn2 = 32'd63; 
32'd2559: dataIn2 = 32'd55; 
32'd2560: dataIn2 = 32'd20; 
32'd2561: dataIn2 = 32'd48; 
32'd2562: dataIn2 = 32'd76; 
32'd2563: dataIn2 = 32'd38; 
32'd2564: dataIn2 = 32'd85; 
32'd2565: dataIn2 = 32'd67; 
32'd2566: dataIn2 = 32'd60; 
32'd2567: dataIn2 = 32'd13; 
32'd2568: dataIn2 = 32'd71; 
32'd2569: dataIn2 = 32'd74; 
32'd2570: dataIn2 = 32'd77; 
32'd2571: dataIn2 = 32'd67; 
32'd2572: dataIn2 = 32'd6; 
32'd2573: dataIn2 = 32'd79; 
32'd2574: dataIn2 = 32'd50; 
32'd2575: dataIn2 = 32'd1; 
32'd2576: dataIn2 = 32'd50; 
32'd2577: dataIn2 = 32'd57; 
32'd2578: dataIn2 = 32'd8; 
32'd2579: dataIn2 = 32'd82; 
32'd2580: dataIn2 = 32'd70; 
32'd2581: dataIn2 = 32'd4; 
32'd2582: dataIn2 = 32'd12; 
32'd2583: dataIn2 = 32'd19; 
32'd2584: dataIn2 = 32'd2; 
32'd2585: dataIn2 = 32'd10; 
32'd2586: dataIn2 = 32'd52; 
32'd2587: dataIn2 = 32'd54; 
32'd2588: dataIn2 = 32'd19; 
32'd2589: dataIn2 = 32'd23; 
32'd2590: dataIn2 = 32'd76; 
32'd2591: dataIn2 = 32'd52; 
32'd2592: dataIn2 = 32'd3; 
32'd2593: dataIn2 = 32'd95; 
32'd2594: dataIn2 = 32'd93; 
32'd2595: dataIn2 = 32'd20; 
32'd2596: dataIn2 = 32'd95; 
32'd2597: dataIn2 = 32'd76; 
32'd2598: dataIn2 = 32'd80; 
32'd2599: dataIn2 = 32'd99; 
32'd2600: dataIn2 = 32'd60; 
32'd2601: dataIn2 = 32'd85; 
32'd2602: dataIn2 = 32'd83; 
32'd2603: dataIn2 = 32'd52; 
32'd2604: dataIn2 = 32'd39; 
32'd2605: dataIn2 = 32'd18; 
32'd2606: dataIn2 = 32'd59; 
32'd2607: dataIn2 = 32'd63; 
32'd2608: dataIn2 = 32'd70; 
32'd2609: dataIn2 = 32'd21; 
32'd2610: dataIn2 = 32'd100; 
32'd2611: dataIn2 = 32'd28; 
32'd2612: dataIn2 = 32'd19; 
32'd2613: dataIn2 = 32'd7; 
32'd2614: dataIn2 = 32'd25; 
32'd2615: dataIn2 = 32'd42; 
32'd2616: dataIn2 = 32'd52; 
32'd2617: dataIn2 = 32'd69; 
32'd2618: dataIn2 = 32'd69; 
32'd2619: dataIn2 = 32'd68; 
32'd2620: dataIn2 = 32'd24; 
32'd2621: dataIn2 = 32'd82; 
32'd2622: dataIn2 = 32'd76; 
32'd2623: dataIn2 = 32'd63; 
32'd2624: dataIn2 = 32'd3; 
32'd2625: dataIn2 = 32'd8; 
32'd2626: dataIn2 = 32'd80; 
32'd2627: dataIn2 = 32'd2; 
32'd2628: dataIn2 = 32'd74; 
32'd2629: dataIn2 = 32'd98; 
32'd2630: dataIn2 = 32'd79; 
32'd2631: dataIn2 = 32'd35; 
32'd2632: dataIn2 = 32'd68; 
32'd2633: dataIn2 = 32'd90; 
32'd2634: dataIn2 = 32'd88; 
32'd2635: dataIn2 = 32'd93; 
32'd2636: dataIn2 = 32'd81; 
32'd2637: dataIn2 = 32'd23; 
32'd2638: dataIn2 = 32'd67; 
32'd2639: dataIn2 = 32'd37; 
32'd2640: dataIn2 = 32'd69; 
32'd2641: dataIn2 = 32'd1; 
32'd2642: dataIn2 = 32'd92; 
32'd2643: dataIn2 = 32'd30; 
32'd2644: dataIn2 = 32'd0; 
32'd2645: dataIn2 = 32'd58; 
32'd2646: dataIn2 = 32'd98; 
32'd2647: dataIn2 = 32'd87; 
32'd2648: dataIn2 = 32'd26; 
32'd2649: dataIn2 = 32'd84; 
32'd2650: dataIn2 = 32'd52; 
32'd2651: dataIn2 = 32'd10; 
32'd2652: dataIn2 = 32'd35; 
32'd2653: dataIn2 = 32'd13; 
32'd2654: dataIn2 = 32'd25; 
32'd2655: dataIn2 = 32'd37; 
32'd2656: dataIn2 = 32'd59; 
32'd2657: dataIn2 = 32'd61; 
32'd2658: dataIn2 = 32'd27; 
32'd2659: dataIn2 = 32'd75; 
32'd2660: dataIn2 = 32'd88; 
32'd2661: dataIn2 = 32'd29; 
32'd2662: dataIn2 = 32'd0; 
32'd2663: dataIn2 = 32'd34; 
32'd2664: dataIn2 = 32'd0; 
32'd2665: dataIn2 = 32'd56; 
32'd2666: dataIn2 = 32'd36; 
32'd2667: dataIn2 = 32'd12; 
32'd2668: dataIn2 = 32'd4; 
32'd2669: dataIn2 = 32'd94; 
32'd2670: dataIn2 = 32'd3; 
32'd2671: dataIn2 = 32'd88; 
32'd2672: dataIn2 = 32'd83; 
32'd2673: dataIn2 = 32'd46; 
32'd2674: dataIn2 = 32'd15; 
32'd2675: dataIn2 = 32'd20; 
32'd2676: dataIn2 = 32'd57; 
32'd2677: dataIn2 = 32'd30; 
32'd2678: dataIn2 = 32'd57; 
32'd2679: dataIn2 = 32'd6; 
32'd2680: dataIn2 = 32'd48; 
32'd2681: dataIn2 = 32'd99; 
32'd2682: dataIn2 = 32'd57; 
32'd2683: dataIn2 = 32'd31; 
32'd2684: dataIn2 = 32'd71; 
32'd2685: dataIn2 = 32'd55; 
32'd2686: dataIn2 = 32'd87; 
32'd2687: dataIn2 = 32'd87; 
32'd2688: dataIn2 = 32'd59; 
32'd2689: dataIn2 = 32'd15; 
32'd2690: dataIn2 = 32'd44; 
32'd2691: dataIn2 = 32'd99; 
32'd2692: dataIn2 = 32'd70; 
32'd2693: dataIn2 = 32'd2; 
32'd2694: dataIn2 = 32'd54; 
32'd2695: dataIn2 = 32'd71; 
32'd2696: dataIn2 = 32'd29; 
32'd2697: dataIn2 = 32'd78; 
32'd2698: dataIn2 = 32'd83; 
32'd2699: dataIn2 = 32'd48; 
32'd2700: dataIn2 = 32'd97; 
32'd2701: dataIn2 = 32'd76; 
32'd2702: dataIn2 = 32'd47; 
32'd2703: dataIn2 = 32'd30; 
32'd2704: dataIn2 = 32'd94; 
32'd2705: dataIn2 = 32'd2; 
32'd2706: dataIn2 = 32'd68; 
32'd2707: dataIn2 = 32'd55; 
32'd2708: dataIn2 = 32'd63; 
32'd2709: dataIn2 = 32'd43; 
32'd2710: dataIn2 = 32'd4; 
32'd2711: dataIn2 = 32'd87; 
32'd2712: dataIn2 = 32'd22; 
32'd2713: dataIn2 = 32'd64; 
32'd2714: dataIn2 = 32'd8; 
32'd2715: dataIn2 = 32'd72; 
32'd2716: dataIn2 = 32'd76; 
32'd2717: dataIn2 = 32'd63; 
32'd2718: dataIn2 = 32'd21; 
32'd2719: dataIn2 = 32'd90; 
32'd2720: dataIn2 = 32'd85; 
32'd2721: dataIn2 = 32'd22; 
32'd2722: dataIn2 = 32'd5; 
32'd2723: dataIn2 = 32'd38; 
32'd2724: dataIn2 = 32'd7; 
32'd2725: dataIn2 = 32'd70; 
32'd2726: dataIn2 = 32'd77; 
32'd2727: dataIn2 = 32'd22; 
32'd2728: dataIn2 = 32'd33; 
32'd2729: dataIn2 = 32'd54; 
32'd2730: dataIn2 = 32'd76; 
32'd2731: dataIn2 = 32'd78; 
32'd2732: dataIn2 = 32'd69; 
32'd2733: dataIn2 = 32'd31; 
32'd2734: dataIn2 = 32'd98; 
32'd2735: dataIn2 = 32'd86; 
32'd2736: dataIn2 = 32'd58; 
32'd2737: dataIn2 = 32'd83; 
32'd2738: dataIn2 = 32'd83; 
32'd2739: dataIn2 = 32'd79; 
32'd2740: dataIn2 = 32'd53; 
32'd2741: dataIn2 = 32'd92; 
32'd2742: dataIn2 = 32'd87; 
32'd2743: dataIn2 = 32'd65; 
32'd2744: dataIn2 = 32'd34; 
32'd2745: dataIn2 = 32'd100; 
32'd2746: dataIn2 = 32'd4; 
32'd2747: dataIn2 = 32'd17; 
32'd2748: dataIn2 = 32'd28; 
32'd2749: dataIn2 = 32'd35; 
32'd2750: dataIn2 = 32'd95; 
32'd2751: dataIn2 = 32'd32; 
32'd2752: dataIn2 = 32'd56; 
32'd2753: dataIn2 = 32'd63; 
32'd2754: dataIn2 = 32'd53; 
32'd2755: dataIn2 = 32'd19; 
32'd2756: dataIn2 = 32'd4; 
32'd2757: dataIn2 = 32'd45; 
32'd2758: dataIn2 = 32'd8; 
32'd2759: dataIn2 = 32'd67; 
32'd2760: dataIn2 = 32'd44; 
32'd2761: dataIn2 = 32'd87; 
32'd2762: dataIn2 = 32'd94; 
32'd2763: dataIn2 = 32'd72; 
32'd2764: dataIn2 = 32'd51; 
32'd2765: dataIn2 = 32'd23; 
32'd2766: dataIn2 = 32'd28; 
32'd2767: dataIn2 = 32'd17; 
32'd2768: dataIn2 = 32'd73; 
32'd2769: dataIn2 = 32'd33; 
32'd2770: dataIn2 = 32'd80; 
32'd2771: dataIn2 = 32'd90; 
32'd2772: dataIn2 = 32'd84; 
32'd2773: dataIn2 = 32'd39; 
32'd2774: dataIn2 = 32'd50; 
32'd2775: dataIn2 = 32'd87; 
32'd2776: dataIn2 = 32'd15; 
32'd2777: dataIn2 = 32'd78; 
32'd2778: dataIn2 = 32'd91; 
32'd2779: dataIn2 = 32'd59; 
32'd2780: dataIn2 = 32'd95; 
32'd2781: dataIn2 = 32'd67; 
32'd2782: dataIn2 = 32'd99; 
32'd2783: dataIn2 = 32'd11; 
32'd2784: dataIn2 = 32'd12; 
32'd2785: dataIn2 = 32'd48; 
32'd2786: dataIn2 = 32'd13; 
32'd2787: dataIn2 = 32'd63; 
32'd2788: dataIn2 = 32'd62; 
32'd2789: dataIn2 = 32'd71; 
32'd2790: dataIn2 = 32'd43; 
32'd2791: dataIn2 = 32'd94; 
32'd2792: dataIn2 = 32'd81; 
32'd2793: dataIn2 = 32'd19; 
32'd2794: dataIn2 = 32'd48; 
32'd2795: dataIn2 = 32'd51; 
32'd2796: dataIn2 = 32'd44; 
32'd2797: dataIn2 = 32'd73; 
32'd2798: dataIn2 = 32'd94; 
32'd2799: dataIn2 = 32'd23; 
32'd2800: dataIn2 = 32'd90; 
32'd2801: dataIn2 = 32'd50; 
32'd2802: dataIn2 = 32'd56; 
32'd2803: dataIn2 = 32'd33; 
32'd2804: dataIn2 = 32'd82; 
32'd2805: dataIn2 = 32'd91; 
32'd2806: dataIn2 = 32'd29; 
32'd2807: dataIn2 = 32'd76; 
32'd2808: dataIn2 = 32'd89; 
32'd2809: dataIn2 = 32'd88; 
32'd2810: dataIn2 = 32'd29; 
32'd2811: dataIn2 = 32'd28; 
32'd2812: dataIn2 = 32'd28; 
32'd2813: dataIn2 = 32'd47; 
32'd2814: dataIn2 = 32'd96; 
32'd2815: dataIn2 = 32'd58; 
32'd2816: dataIn2 = 32'd100; 
32'd2817: dataIn2 = 32'd16; 
32'd2818: dataIn2 = 32'd14; 
32'd2819: dataIn2 = 32'd46; 
32'd2820: dataIn2 = 32'd60; 
32'd2821: dataIn2 = 32'd4; 
32'd2822: dataIn2 = 32'd53; 
32'd2823: dataIn2 = 32'd59; 
32'd2824: dataIn2 = 32'd0; 
32'd2825: dataIn2 = 32'd98; 
32'd2826: dataIn2 = 32'd54; 
32'd2827: dataIn2 = 32'd60; 
32'd2828: dataIn2 = 32'd81; 
32'd2829: dataIn2 = 32'd40; 
32'd2830: dataIn2 = 32'd54; 
32'd2831: dataIn2 = 32'd59; 
32'd2832: dataIn2 = 32'd8; 
32'd2833: dataIn2 = 32'd0; 
32'd2834: dataIn2 = 32'd55; 
32'd2835: dataIn2 = 32'd87; 
32'd2836: dataIn2 = 32'd87; 
32'd2837: dataIn2 = 32'd15; 
32'd2838: dataIn2 = 32'd21; 
32'd2839: dataIn2 = 32'd6; 
32'd2840: dataIn2 = 32'd80; 
32'd2841: dataIn2 = 32'd46; 
32'd2842: dataIn2 = 32'd40; 
32'd2843: dataIn2 = 32'd87; 
32'd2844: dataIn2 = 32'd18; 
32'd2845: dataIn2 = 32'd13; 
32'd2846: dataIn2 = 32'd10; 
32'd2847: dataIn2 = 32'd50; 
32'd2848: dataIn2 = 32'd10; 
32'd2849: dataIn2 = 32'd57; 
32'd2850: dataIn2 = 32'd96; 
32'd2851: dataIn2 = 32'd43; 
32'd2852: dataIn2 = 32'd14; 
32'd2853: dataIn2 = 32'd68; 
32'd2854: dataIn2 = 32'd85; 
32'd2855: dataIn2 = 32'd24; 
32'd2856: dataIn2 = 32'd26; 
32'd2857: dataIn2 = 32'd29; 
32'd2858: dataIn2 = 32'd41; 
32'd2859: dataIn2 = 32'd40; 
32'd2860: dataIn2 = 32'd58; 
32'd2861: dataIn2 = 32'd23; 
32'd2862: dataIn2 = 32'd13; 
32'd2863: dataIn2 = 32'd17; 
32'd2864: dataIn2 = 32'd17; 
32'd2865: dataIn2 = 32'd67; 
32'd2866: dataIn2 = 32'd26; 
32'd2867: dataIn2 = 32'd60; 
32'd2868: dataIn2 = 32'd43; 
32'd2869: dataIn2 = 32'd9; 
32'd2870: dataIn2 = 32'd39; 
32'd2871: dataIn2 = 32'd80; 
32'd2872: dataIn2 = 32'd43; 
32'd2873: dataIn2 = 32'd82; 
32'd2874: dataIn2 = 32'd88; 
32'd2875: dataIn2 = 32'd21; 
32'd2876: dataIn2 = 32'd87; 
32'd2877: dataIn2 = 32'd25; 
32'd2878: dataIn2 = 32'd54; 
32'd2879: dataIn2 = 32'd78; 
32'd2880: dataIn2 = 32'd51; 
32'd2881: dataIn2 = 32'd97; 
32'd2882: dataIn2 = 32'd13; 
32'd2883: dataIn2 = 32'd73; 
32'd2884: dataIn2 = 32'd35; 
32'd2885: dataIn2 = 32'd94; 
32'd2886: dataIn2 = 32'd68; 
32'd2887: dataIn2 = 32'd57; 
32'd2888: dataIn2 = 32'd59; 
32'd2889: dataIn2 = 32'd77; 
32'd2890: dataIn2 = 32'd5; 
32'd2891: dataIn2 = 32'd79; 
32'd2892: dataIn2 = 32'd28; 
32'd2893: dataIn2 = 32'd68; 
32'd2894: dataIn2 = 32'd93; 
32'd2895: dataIn2 = 32'd99; 
32'd2896: dataIn2 = 32'd70; 
32'd2897: dataIn2 = 32'd67; 
32'd2898: dataIn2 = 32'd18; 
32'd2899: dataIn2 = 32'd32; 
32'd2900: dataIn2 = 32'd41; 
32'd2901: dataIn2 = 32'd62; 
32'd2902: dataIn2 = 32'd67; 
32'd2903: dataIn2 = 32'd91; 
32'd2904: dataIn2 = 32'd54; 
32'd2905: dataIn2 = 32'd86; 
32'd2906: dataIn2 = 32'd71; 
32'd2907: dataIn2 = 32'd39; 
32'd2908: dataIn2 = 32'd25; 
32'd2909: dataIn2 = 32'd69; 
32'd2910: dataIn2 = 32'd15; 
32'd2911: dataIn2 = 32'd50; 
32'd2912: dataIn2 = 32'd39; 
32'd2913: dataIn2 = 32'd23; 
32'd2914: dataIn2 = 32'd84; 
32'd2915: dataIn2 = 32'd69; 
32'd2916: dataIn2 = 32'd1; 
32'd2917: dataIn2 = 32'd6; 
32'd2918: dataIn2 = 32'd6; 
32'd2919: dataIn2 = 32'd16; 
32'd2920: dataIn2 = 32'd57; 
32'd2921: dataIn2 = 32'd98; 
32'd2922: dataIn2 = 32'd17; 
32'd2923: dataIn2 = 32'd36; 
32'd2924: dataIn2 = 32'd8; 
32'd2925: dataIn2 = 32'd95; 
32'd2926: dataIn2 = 32'd69; 
32'd2927: dataIn2 = 32'd12; 
32'd2928: dataIn2 = 32'd37; 
32'd2929: dataIn2 = 32'd77; 
32'd2930: dataIn2 = 32'd89; 
32'd2931: dataIn2 = 32'd77; 
32'd2932: dataIn2 = 32'd28; 
32'd2933: dataIn2 = 32'd29; 
32'd2934: dataIn2 = 32'd36; 
32'd2935: dataIn2 = 32'd26; 
32'd2936: dataIn2 = 32'd34; 
32'd2937: dataIn2 = 32'd86; 
32'd2938: dataIn2 = 32'd65; 
32'd2939: dataIn2 = 32'd61; 
32'd2940: dataIn2 = 32'd74; 
32'd2941: dataIn2 = 32'd27; 
32'd2942: dataIn2 = 32'd75; 
32'd2943: dataIn2 = 32'd67; 
32'd2944: dataIn2 = 32'd37; 
32'd2945: dataIn2 = 32'd31; 
32'd2946: dataIn2 = 32'd41; 
32'd2947: dataIn2 = 32'd68; 
32'd2948: dataIn2 = 32'd29; 
32'd2949: dataIn2 = 32'd46; 
32'd2950: dataIn2 = 32'd63; 
32'd2951: dataIn2 = 32'd46; 
32'd2952: dataIn2 = 32'd86; 
32'd2953: dataIn2 = 32'd33; 
32'd2954: dataIn2 = 32'd3; 
32'd2955: dataIn2 = 32'd97; 
32'd2956: dataIn2 = 32'd86; 
32'd2957: dataIn2 = 32'd50; 
32'd2958: dataIn2 = 32'd88; 
32'd2959: dataIn2 = 32'd23; 
32'd2960: dataIn2 = 32'd82; 
32'd2961: dataIn2 = 32'd92; 
32'd2962: dataIn2 = 32'd79; 
32'd2963: dataIn2 = 32'd91; 
32'd2964: dataIn2 = 32'd52; 
32'd2965: dataIn2 = 32'd44; 
32'd2966: dataIn2 = 32'd87; 
32'd2967: dataIn2 = 32'd54; 
32'd2968: dataIn2 = 32'd90; 
32'd2969: dataIn2 = 32'd38; 
32'd2970: dataIn2 = 32'd0; 
32'd2971: dataIn2 = 32'd27; 
32'd2972: dataIn2 = 32'd93; 
32'd2973: dataIn2 = 32'd52; 
32'd2974: dataIn2 = 32'd34; 
32'd2975: dataIn2 = 32'd16; 
32'd2976: dataIn2 = 32'd76; 
32'd2977: dataIn2 = 32'd28; 
32'd2978: dataIn2 = 32'd95; 
32'd2979: dataIn2 = 32'd27; 
32'd2980: dataIn2 = 32'd72; 
32'd2981: dataIn2 = 32'd84; 
32'd2982: dataIn2 = 32'd93; 
32'd2983: dataIn2 = 32'd23; 
32'd2984: dataIn2 = 32'd20; 
32'd2985: dataIn2 = 32'd82; 
32'd2986: dataIn2 = 32'd84; 
32'd2987: dataIn2 = 32'd64; 
32'd2988: dataIn2 = 32'd80; 
32'd2989: dataIn2 = 32'd29; 
32'd2990: dataIn2 = 32'd77; 
32'd2991: dataIn2 = 32'd99; 
32'd2992: dataIn2 = 32'd9; 
32'd2993: dataIn2 = 32'd70; 
32'd2994: dataIn2 = 32'd83; 
32'd2995: dataIn2 = 32'd91; 
32'd2996: dataIn2 = 32'd28; 
32'd2997: dataIn2 = 32'd51; 
32'd2998: dataIn2 = 32'd78; 
32'd2999: dataIn2 = 32'd57; 
32'd3000: dataIn2 = 32'd41; 
32'd3001: dataIn2 = 32'd4; 
32'd3002: dataIn2 = 32'd29; 
32'd3003: dataIn2 = 32'd1; 
32'd3004: dataIn2 = 32'd22; 
32'd3005: dataIn2 = 32'd18; 
32'd3006: dataIn2 = 32'd80; 
32'd3007: dataIn2 = 32'd96; 
32'd3008: dataIn2 = 32'd29; 
32'd3009: dataIn2 = 32'd48; 
32'd3010: dataIn2 = 32'd36; 
32'd3011: dataIn2 = 32'd14; 
32'd3012: dataIn2 = 32'd26; 
32'd3013: dataIn2 = 32'd88; 
32'd3014: dataIn2 = 32'd64; 
32'd3015: dataIn2 = 32'd50; 
32'd3016: dataIn2 = 32'd20; 
32'd3017: dataIn2 = 32'd91; 
32'd3018: dataIn2 = 32'd38; 
32'd3019: dataIn2 = 32'd63; 
32'd3020: dataIn2 = 32'd19; 
32'd3021: dataIn2 = 32'd94; 
32'd3022: dataIn2 = 32'd69; 
32'd3023: dataIn2 = 32'd90; 
32'd3024: dataIn2 = 32'd44; 
32'd3025: dataIn2 = 32'd42; 
32'd3026: dataIn2 = 32'd8; 
32'd3027: dataIn2 = 32'd48; 
32'd3028: dataIn2 = 32'd92; 
32'd3029: dataIn2 = 32'd13; 
32'd3030: dataIn2 = 32'd86; 
32'd3031: dataIn2 = 32'd50; 
32'd3032: dataIn2 = 32'd45; 
32'd3033: dataIn2 = 32'd87; 
32'd3034: dataIn2 = 32'd36; 
32'd3035: dataIn2 = 32'd82; 
32'd3036: dataIn2 = 32'd15; 
32'd3037: dataIn2 = 32'd75; 
32'd3038: dataIn2 = 32'd41; 
32'd3039: dataIn2 = 32'd82; 
32'd3040: dataIn2 = 32'd13; 
32'd3041: dataIn2 = 32'd67; 
32'd3042: dataIn2 = 32'd17; 
32'd3043: dataIn2 = 32'd16; 
32'd3044: dataIn2 = 32'd98; 
32'd3045: dataIn2 = 32'd53; 
32'd3046: dataIn2 = 32'd8; 
32'd3047: dataIn2 = 32'd2; 
32'd3048: dataIn2 = 32'd89; 
32'd3049: dataIn2 = 32'd16; 
32'd3050: dataIn2 = 32'd0; 
32'd3051: dataIn2 = 32'd33; 
32'd3052: dataIn2 = 32'd81; 
32'd3053: dataIn2 = 32'd28; 
32'd3054: dataIn2 = 32'd92; 
32'd3055: dataIn2 = 32'd76; 
32'd3056: dataIn2 = 32'd66; 
32'd3057: dataIn2 = 32'd72; 
32'd3058: dataIn2 = 32'd98; 
32'd3059: dataIn2 = 32'd38; 
32'd3060: dataIn2 = 32'd71; 
32'd3061: dataIn2 = 32'd63; 
32'd3062: dataIn2 = 32'd57; 
32'd3063: dataIn2 = 32'd83; 
32'd3064: dataIn2 = 32'd17; 
32'd3065: dataIn2 = 32'd94; 
32'd3066: dataIn2 = 32'd89; 
32'd3067: dataIn2 = 32'd33; 
32'd3068: dataIn2 = 32'd43; 
32'd3069: dataIn2 = 32'd87; 
32'd3070: dataIn2 = 32'd91; 
32'd3071: dataIn2 = 32'd15; 
32'd3072: dataIn2 = 32'd38; 
32'd3073: dataIn2 = 32'd93; 
32'd3074: dataIn2 = 32'd23; 
32'd3075: dataIn2 = 32'd49; 
32'd3076: dataIn2 = 32'd16; 
32'd3077: dataIn2 = 32'd66; 
32'd3078: dataIn2 = 32'd65; 
32'd3079: dataIn2 = 32'd62; 
32'd3080: dataIn2 = 32'd53; 
32'd3081: dataIn2 = 32'd75; 
32'd3082: dataIn2 = 32'd9; 
32'd3083: dataIn2 = 32'd78; 
32'd3084: dataIn2 = 32'd35; 
32'd3085: dataIn2 = 32'd5; 
32'd3086: dataIn2 = 32'd23; 
32'd3087: dataIn2 = 32'd66; 
32'd3088: dataIn2 = 32'd86; 
32'd3089: dataIn2 = 32'd74; 
32'd3090: dataIn2 = 32'd72; 
32'd3091: dataIn2 = 32'd36; 
32'd3092: dataIn2 = 32'd7; 
32'd3093: dataIn2 = 32'd29; 
32'd3094: dataIn2 = 32'd29; 
32'd3095: dataIn2 = 32'd44; 
32'd3096: dataIn2 = 32'd80; 
32'd3097: dataIn2 = 32'd80; 
32'd3098: dataIn2 = 32'd6; 
32'd3099: dataIn2 = 32'd11; 
32'd3100: dataIn2 = 32'd13; 
32'd3101: dataIn2 = 32'd71; 
32'd3102: dataIn2 = 32'd14; 
32'd3103: dataIn2 = 32'd90; 
32'd3104: dataIn2 = 32'd53; 
32'd3105: dataIn2 = 32'd77; 
32'd3106: dataIn2 = 32'd81; 
32'd3107: dataIn2 = 32'd85; 
32'd3108: dataIn2 = 32'd59; 
32'd3109: dataIn2 = 32'd20; 
32'd3110: dataIn2 = 32'd29; 
32'd3111: dataIn2 = 32'd77; 
32'd3112: dataIn2 = 32'd61; 
32'd3113: dataIn2 = 32'd49; 
32'd3114: dataIn2 = 32'd74; 
32'd3115: dataIn2 = 32'd89; 
32'd3116: dataIn2 = 32'd54; 
32'd3117: dataIn2 = 32'd34; 
32'd3118: dataIn2 = 32'd5; 
32'd3119: dataIn2 = 32'd75; 
32'd3120: dataIn2 = 32'd76; 
32'd3121: dataIn2 = 32'd48; 
32'd3122: dataIn2 = 32'd22; 
32'd3123: dataIn2 = 32'd53; 
32'd3124: dataIn2 = 32'd97; 
32'd3125: dataIn2 = 32'd28; 
32'd3126: dataIn2 = 32'd81; 
32'd3127: dataIn2 = 32'd19; 
32'd3128: dataIn2 = 32'd96; 
32'd3129: dataIn2 = 32'd54; 
32'd3130: dataIn2 = 32'd8; 
32'd3131: dataIn2 = 32'd79; 
32'd3132: dataIn2 = 32'd15; 
32'd3133: dataIn2 = 32'd52; 
32'd3134: dataIn2 = 32'd45; 
32'd3135: dataIn2 = 32'd30; 
32'd3136: dataIn2 = 32'd11; 
32'd3137: dataIn2 = 32'd91; 
32'd3138: dataIn2 = 32'd20; 
32'd3139: dataIn2 = 32'd51; 
32'd3140: dataIn2 = 32'd67; 
32'd3141: dataIn2 = 32'd92; 
32'd3142: dataIn2 = 32'd31; 
32'd3143: dataIn2 = 32'd21; 
32'd3144: dataIn2 = 32'd57; 
32'd3145: dataIn2 = 32'd18; 
32'd3146: dataIn2 = 32'd74; 
32'd3147: dataIn2 = 32'd23; 
32'd3148: dataIn2 = 32'd26; 
32'd3149: dataIn2 = 32'd50; 
32'd3150: dataIn2 = 32'd58; 
32'd3151: dataIn2 = 32'd16; 
32'd3152: dataIn2 = 32'd65; 
32'd3153: dataIn2 = 32'd15; 
32'd3154: dataIn2 = 32'd86; 
32'd3155: dataIn2 = 32'd49; 
32'd3156: dataIn2 = 32'd30; 
32'd3157: dataIn2 = 32'd21; 
32'd3158: dataIn2 = 32'd13; 
32'd3159: dataIn2 = 32'd34; 
32'd3160: dataIn2 = 32'd42; 
32'd3161: dataIn2 = 32'd76; 
32'd3162: dataIn2 = 32'd33; 
32'd3163: dataIn2 = 32'd10; 
32'd3164: dataIn2 = 32'd90; 
32'd3165: dataIn2 = 32'd63; 
32'd3166: dataIn2 = 32'd15; 
32'd3167: dataIn2 = 32'd36; 
32'd3168: dataIn2 = 32'd33; 
32'd3169: dataIn2 = 32'd88; 
32'd3170: dataIn2 = 32'd99; 
32'd3171: dataIn2 = 32'd76; 
32'd3172: dataIn2 = 32'd54; 
32'd3173: dataIn2 = 32'd53; 
32'd3174: dataIn2 = 32'd7; 
32'd3175: dataIn2 = 32'd53; 
32'd3176: dataIn2 = 32'd94; 
32'd3177: dataIn2 = 32'd40; 
32'd3178: dataIn2 = 32'd85; 
32'd3179: dataIn2 = 32'd20; 
32'd3180: dataIn2 = 32'd18; 
32'd3181: dataIn2 = 32'd33; 
32'd3182: dataIn2 = 32'd70; 
32'd3183: dataIn2 = 32'd6; 
32'd3184: dataIn2 = 32'd1; 
32'd3185: dataIn2 = 32'd11; 
32'd3186: dataIn2 = 32'd52; 
32'd3187: dataIn2 = 32'd65; 
32'd3188: dataIn2 = 32'd72; 
32'd3189: dataIn2 = 32'd95; 
32'd3190: dataIn2 = 32'd71; 
32'd3191: dataIn2 = 32'd83; 
32'd3192: dataIn2 = 32'd27; 
32'd3193: dataIn2 = 32'd96; 
32'd3194: dataIn2 = 32'd50; 
32'd3195: dataIn2 = 32'd75; 
32'd3196: dataIn2 = 32'd75; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_64_30.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
