//32x32 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 717 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,addr1,addr2,dataIn1,dataIn2,Rst,csize,RD);  
//frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  wdata_col_base = 32'd340 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #122000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd340: dataIn1 = 32'd7; 
32'd341: dataIn1 = 32'd20; 
32'd342: dataIn1 = 32'd1; 
32'd343: dataIn1 = 32'd21; 
32'd344: dataIn1 = 32'd25; 
32'd345: dataIn1 = 32'd7; 
32'd346: dataIn1 = 32'd14; 
32'd347: dataIn1 = 32'd26; 
32'd348: dataIn1 = 32'd4; 
32'd349: dataIn1 = 32'd10; 
32'd350: dataIn1 = 32'd11; 
32'd351: dataIn1 = 32'd25; 
32'd352: dataIn1 = 32'd8; 
32'd353: dataIn1 = 32'd22; 
32'd354: dataIn1 = 32'd15; 
32'd355: dataIn1 = 32'd9; 
32'd356: dataIn1 = 32'd20; 
32'd357: dataIn1 = 32'd12; 
32'd358: dataIn1 = 32'd27; 
32'd359: dataIn1 = 32'd25; 
32'd360: dataIn1 = 32'd24; 
32'd361: dataIn1 = 32'd4; 
32'd362: dataIn1 = 32'd24; 
32'd363: dataIn1 = 32'd2; 
32'd364: dataIn1 = 32'd25; 
32'd365: dataIn1 = 32'd11; 
32'd366: dataIn1 = 32'd5; 
32'd367: dataIn1 = 32'd4; 
32'd368: dataIn1 = 32'd2; 
32'd369: dataIn1 = 32'd21; 
32'd370: dataIn1 = 32'd30; 
32'd371: dataIn1 = 32'd19; 
32'd372: dataIn1 = 32'd29; 
32'd373: dataIn1 = 32'd12; 
32'd374: dataIn1 = 32'd18; 
32'd375: dataIn1 = 32'd27; 
32'd376: dataIn1 = 32'd20; 
32'd377: dataIn1 = 32'd8; 
32'd378: dataIn1 = 32'd16; 
32'd379: dataIn1 = 32'd14; 
32'd380: dataIn1 = 32'd25; 
32'd381: dataIn1 = 32'd13; 
32'd382: dataIn1 = 32'd1; 
32'd383: dataIn1 = 32'd13; 
32'd384: dataIn1 = 32'd9; 
32'd385: dataIn1 = 32'd19; 
32'd386: dataIn1 = 32'd18; 
32'd387: dataIn1 = 32'd22; 
32'd388: dataIn1 = 32'd9; 
32'd389: dataIn1 = 32'd16; 
32'd390: dataIn1 = 32'd1; 
32'd391: dataIn1 = 32'd19; 
32'd392: dataIn1 = 32'd23; 
32'd393: dataIn1 = 32'd3; 
32'd394: dataIn1 = 32'd1; 
32'd395: dataIn1 = 32'd11; 
32'd396: dataIn1 = 32'd13; 
32'd397: dataIn1 = 32'd7; 
32'd398: dataIn1 = 32'd2; 
32'd399: dataIn1 = 32'd10; 
32'd400: dataIn1 = 32'd15; 
32'd401: dataIn1 = 32'd7; 
32'd402: dataIn1 = 32'd6; 
32'd403: dataIn1 = 32'd27; 
32'd404: dataIn1 = 32'd27; 
32'd405: dataIn1 = 32'd4; 
32'd406: dataIn1 = 32'd16; 
32'd407: dataIn1 = 32'd16; 
32'd408: dataIn1 = 32'd1; 
32'd409: dataIn1 = 32'd30; 
32'd410: dataIn1 = 32'd26; 
32'd411: dataIn1 = 32'd11; 
32'd412: dataIn1 = 32'd9; 
32'd413: dataIn1 = 32'd21; 
32'd414: dataIn1 = 32'd3; 
32'd415: dataIn1 = 32'd28; 
32'd416: dataIn1 = 32'd19; 
32'd417: dataIn1 = 32'd24; 
32'd418: dataIn1 = 32'd27; 
32'd419: dataIn1 = 32'd9; 
32'd420: dataIn1 = 32'd28; 
32'd421: dataIn1 = 32'd1; 
32'd422: dataIn1 = 32'd8; 
32'd423: dataIn1 = 32'd11; 
32'd424: dataIn1 = 32'd7; 
32'd425: dataIn1 = 32'd31; 
32'd426: dataIn1 = 32'd25; 
32'd427: dataIn1 = 32'd6; 
32'd428: dataIn1 = 32'd2; 
32'd429: dataIn1 = 32'd14; 
32'd430: dataIn1 = 32'd0; 
32'd431: dataIn1 = 32'd17; 
32'd432: dataIn1 = 32'd24; 
32'd433: dataIn1 = 32'd31; 
32'd434: dataIn1 = 32'd1; 
32'd435: dataIn1 = 32'd14; 
32'd436: dataIn1 = 32'd9; 
32'd437: dataIn1 = 32'd22; 
32'd438: dataIn1 = 32'd0; 
32'd439: dataIn1 = 32'd6; 
32'd440: dataIn1 = 32'd13; 
32'd441: dataIn1 = 32'd13; 
32'd442: dataIn1 = 32'd9; 
32'd443: dataIn1 = 32'd0; 
32'd444: dataIn1 = 32'd14; 
32'd445: dataIn1 = 32'd14; 
32'd446: dataIn1 = 32'd25; 
32'd447: dataIn1 = 32'd10; 
32'd448: dataIn1 = 32'd8; 
32'd449: dataIn1 = 32'd12; 
32'd450: dataIn1 = 32'd5; 
32'd451: dataIn1 = 32'd11; 
32'd452: dataIn1 = 32'd31; 
32'd453: dataIn1 = 32'd8; 
32'd454: dataIn1 = 32'd10; 
32'd455: dataIn1 = 32'd27; 
32'd456: dataIn1 = 32'd31; 
32'd457: dataIn1 = 32'd3; 
32'd458: dataIn1 = 32'd25; 
32'd459: dataIn1 = 32'd30; 
32'd460: dataIn1 = 32'd18; 
32'd461: dataIn1 = 32'd22; 
32'd462: dataIn1 = 32'd1; 
32'd463: dataIn1 = 32'd16; 
32'd464: dataIn1 = 32'd11; 
32'd465: dataIn1 = 32'd7; 
32'd466: dataIn1 = 32'd9; 
32'd467: dataIn1 = 32'd25; 
32'd468: dataIn1 = 32'd27; 
32'd469: dataIn1 = 32'd31; 
32'd470: dataIn1 = 32'd0; 
32'd471: dataIn1 = 32'd20; 
32'd472: dataIn1 = 32'd20; 
32'd473: dataIn1 = 32'd19; 
32'd474: dataIn1 = 32'd21; 
32'd475: dataIn1 = 32'd27; 
32'd476: dataIn1 = 32'd0; 
32'd477: dataIn1 = 32'd25; 
32'd478: dataIn1 = 32'd28; 
32'd479: dataIn1 = 32'd29; 
32'd480: dataIn1 = 32'd13; 
32'd481: dataIn1 = 32'd21; 
32'd482: dataIn1 = 32'd3; 
32'd483: dataIn1 = 32'd5; 
32'd484: dataIn1 = 32'd9; 
32'd485: dataIn1 = 32'd5; 
32'd486: dataIn1 = 32'd4; 
32'd487: dataIn1 = 32'd30; 
32'd488: dataIn1 = 32'd28; 
32'd489: dataIn1 = 32'd1; 
32'd490: dataIn1 = 32'd18; 
32'd491: dataIn1 = 32'd0; 
32'd492: dataIn1 = 32'd11; 
32'd493: dataIn1 = 32'd9; 
32'd494: dataIn1 = 32'd4; 
32'd495: dataIn1 = 32'd17; 
32'd496: dataIn1 = 32'd4; 
32'd497: dataIn1 = 32'd30; 
32'd498: dataIn1 = 32'd30; 
32'd499: dataIn1 = 32'd9; 
32'd500: dataIn1 = 32'd12; 
32'd501: dataIn1 = 32'd22; 
32'd502: dataIn1 = 32'd18; 
32'd503: dataIn1 = 32'd2; 
32'd504: dataIn1 = 32'd28; 
32'd505: dataIn1 = 32'd1; 
32'd506: dataIn1 = 32'd5; 
32'd507: dataIn1 = 32'd6; 
32'd508: dataIn1 = 32'd11; 
32'd509: dataIn1 = 32'd21; 
32'd510: dataIn1 = 32'd18; 
32'd511: dataIn1 = 32'd19; 
32'd512: dataIn1 = 32'd11; 
32'd513: dataIn1 = 32'd29; 
32'd514: dataIn1 = 32'd19; 
32'd515: dataIn1 = 32'd9; 
32'd516: dataIn1 = 32'd17; 
32'd517: dataIn1 = 32'd15; 
32'd518: dataIn1 = 32'd1; 
32'd519: dataIn1 = 32'd6; 
32'd520: dataIn1 = 32'd3; 
32'd521: dataIn1 = 32'd31; 
32'd522: dataIn1 = 32'd7; 
32'd523: dataIn1 = 32'd18; 
32'd524: dataIn1 = 32'd9; 
32'd525: dataIn1 = 32'd25; 
32'd526: dataIn1 = 32'd18; 
32'd527: dataIn1 = 32'd17; 
32'd528: dataIn1 = 32'd14; 
32'd529: dataIn1 = 32'd18; 
32'd530: dataIn1 = 32'd12; 
32'd531: dataIn1 = 32'd30; 
32'd532: dataIn1 = 32'd27; 
32'd533: dataIn1 = 32'd2; 
32'd534: dataIn1 = 32'd26; 
32'd535: dataIn1 = 32'd27; 
32'd536: dataIn1 = 32'd0; 
32'd537: dataIn1 = 32'd23; 
32'd538: dataIn1 = 32'd20; 
32'd539: dataIn1 = 32'd30; 
32'd540: dataIn1 = 32'd17; 
32'd541: dataIn1 = 32'd16; 
32'd542: dataIn1 = 32'd21; 
32'd543: dataIn1 = 32'd8; 
32'd544: dataIn1 = 32'd1; 
32'd545: dataIn1 = 32'd29; 
32'd546: dataIn1 = 32'd8; 
32'd547: dataIn1 = 32'd3; 
32'd548: dataIn1 = 32'd5; 
32'd549: dataIn1 = 32'd11; 
32'd550: dataIn1 = 32'd17; 
32'd551: dataIn1 = 32'd24; 
32'd552: dataIn1 = 32'd5; 
32'd553: dataIn1 = 32'd4; 
32'd554: dataIn1 = 32'd31; 
32'd555: dataIn1 = 32'd5; 
32'd556: dataIn1 = 32'd30; 
32'd557: dataIn1 = 32'd12; 
32'd558: dataIn1 = 32'd16; 
32'd559: dataIn1 = 32'd13; 
32'd560: dataIn1 = 32'd12; 
32'd561: dataIn1 = 32'd0; 
32'd562: dataIn1 = 32'd6; 
32'd563: dataIn1 = 32'd1; 
32'd564: dataIn1 = 32'd14; 
32'd565: dataIn1 = 32'd22; 
32'd566: dataIn1 = 32'd5; 
32'd567: dataIn1 = 32'd10; 
32'd568: dataIn1 = 32'd27; 
32'd569: dataIn1 = 32'd3; 
32'd570: dataIn1 = 32'd12; 
32'd571: dataIn1 = 32'd0; 
32'd572: dataIn1 = 32'd5; 
32'd573: dataIn1 = 32'd31; 
32'd574: dataIn1 = 32'd13; 
32'd575: dataIn1 = 32'd31; 
32'd576: dataIn1 = 32'd16; 
32'd577: dataIn1 = 32'd21; 
32'd578: dataIn1 = 32'd2; 
32'd579: dataIn1 = 32'd0; 
32'd580: dataIn1 = 32'd21; 
32'd581: dataIn1 = 32'd16; 
32'd582: dataIn1 = 32'd0; 
32'd583: dataIn1 = 32'd6; 
32'd584: dataIn1 = 32'd18; 
32'd585: dataIn1 = 32'd26; 
32'd586: dataIn1 = 32'd3; 
32'd587: dataIn1 = 32'd1; 
32'd588: dataIn1 = 32'd4; 
32'd589: dataIn1 = 32'd3; 
32'd590: dataIn1 = 32'd20; 
32'd591: dataIn1 = 32'd26; 
32'd592: dataIn1 = 32'd4; 
32'd593: dataIn1 = 32'd15; 
32'd594: dataIn1 = 32'd26; 
32'd595: dataIn1 = 32'd6; 
32'd596: dataIn1 = 32'd20; 
32'd597: dataIn1 = 32'd5; 
32'd598: dataIn1 = 32'd1; 
32'd599: dataIn1 = 32'd9; 
32'd600: dataIn1 = 32'd29; 
32'd601: dataIn1 = 32'd25; 
32'd602: dataIn1 = 32'd30; 
32'd603: dataIn1 = 32'd10; 
32'd604: dataIn1 = 32'd14; 
32'd605: dataIn1 = 32'd7; 
32'd606: dataIn1 = 32'd0; 
32'd607: dataIn1 = 32'd4; 
32'd608: dataIn1 = 32'd4; 
32'd609: dataIn1 = 32'd12; 
32'd610: dataIn1 = 32'd30; 
32'd611: dataIn1 = 32'd23; 
32'd612: dataIn1 = 32'd31; 
32'd613: dataIn1 = 32'd7; 
32'd614: dataIn1 = 32'd29; 
32'd615: dataIn1 = 32'd12; 
32'd616: dataIn1 = 32'd12; 
32'd617: dataIn1 = 32'd1; 
32'd618: dataIn1 = 32'd11; 
32'd619: dataIn1 = 32'd25; 
32'd620: dataIn1 = 32'd4; 
32'd621: dataIn1 = 32'd27; 
32'd622: dataIn1 = 32'd4; 
32'd623: dataIn1 = 32'd10; 
32'd624: dataIn1 = 32'd30; 
32'd625: dataIn1 = 32'd26; 
32'd626: dataIn1 = 32'd14; 
32'd627: dataIn1 = 32'd13; 
32'd628: dataIn1 = 32'd6; 
32'd629: dataIn1 = 32'd17; 
32'd630: dataIn1 = 32'd2; 
32'd631: dataIn1 = 32'd9; 
32'd632: dataIn1 = 32'd18; 
32'd633: dataIn1 = 32'd20; 
32'd634: dataIn1 = 32'd27; 
32'd635: dataIn1 = 32'd29; 
32'd636: dataIn1 = 32'd0; 
32'd637: dataIn1 = 32'd20; 
32'd638: dataIn1 = 32'd29; 
32'd639: dataIn1 = 32'd13; 
32'd640: dataIn1 = 32'd0; 
32'd641: dataIn1 = 32'd11; 
32'd642: dataIn1 = 32'd8; 
32'd643: dataIn1 = 32'd10; 
32'd644: dataIn1 = 32'd27; 
32'd645: dataIn1 = 32'd4; 
32'd646: dataIn1 = 32'd19; 
32'd647: dataIn1 = 32'd12; 
32'd648: dataIn1 = 32'd22; 
32'd649: dataIn1 = 32'd29; 
32'd650: dataIn1 = 32'd13; 
32'd651: dataIn1 = 32'd10; 
32'd652: dataIn1 = 32'd24; 
32'd653: dataIn1 = 32'd20; 
32'd654: dataIn1 = 32'd5; 
32'd655: dataIn1 = 32'd11; 
32'd656: dataIn1 = 32'd26; 
32'd657: dataIn1 = 32'd28; 
32'd658: dataIn1 = 32'd4; 
32'd659: dataIn1 = 32'd18; 
32'd660: dataIn1 = 32'd2; 
32'd661: dataIn1 = 32'd21; 
32'd662: dataIn1 = 32'd27; 
32'd663: dataIn1 = 32'd11; 
32'd664: dataIn1 = 32'd20; 
32'd665: dataIn1 = 32'd30; 
32'd666: dataIn1 = 32'd7; 
32'd667: dataIn1 = 32'd19; 
32'd668: dataIn1 = 32'd5; 
32'd669: dataIn1 = 32'd15; 
32'd670: dataIn1 = 32'd3; 
32'd671: dataIn1 = 32'd5; 
32'd672: dataIn1 = 32'd20; 
32'd673: dataIn1 = 32'd31; 
32'd674: dataIn1 = 32'd13; 
32'd675: dataIn1 = 32'd17; 
32'd676: dataIn1 = 32'd2; 
32'd677: dataIn1 = 32'd23; 
32'd678: dataIn1 = 32'd21; 
32'd679: dataIn1 = 32'd18; 
32'd680: dataIn1 = 32'd17; 
32'd681: dataIn1 = 32'd17; 
32'd682: dataIn1 = 32'd7; 
32'd683: dataIn1 = 32'd7; 
32'd684: dataIn1 = 32'd29; 
32'd685: dataIn1 = 32'd24; 
32'd686: dataIn1 = 32'd22; 
32'd687: dataIn1 = 32'd31; 
32'd688: dataIn1 = 32'd21; 
32'd689: dataIn1 = 32'd0; 
32'd690: dataIn1 = 32'd18; 
32'd691: dataIn1 = 32'd4; 
32'd692: dataIn1 = 32'd25; 
32'd693: dataIn1 = 32'd22; 
32'd694: dataIn1 = 32'd16; 
32'd695: dataIn1 = 32'd31; 
32'd696: dataIn1 = 32'd21; 
32'd697: dataIn1 = 32'd18; 
32'd698: dataIn1 = 32'd31; 
32'd699: dataIn1 = 32'd0; 
32'd700: dataIn1 = 32'd30; 
32'd701: dataIn1 = 32'd15; 
32'd702: dataIn1 = 32'd10; 
32'd703: dataIn1 = 32'd11; 
32'd704: dataIn1 = 32'd21; 
32'd705: dataIn1 = 32'd11; 
32'd706: dataIn1 = 32'd30; 
32'd707: dataIn1 = 32'd18; 
32'd708: dataIn1 = 32'd20; 
32'd709: dataIn1 = 32'd28; 
32'd710: dataIn1 = 32'd30; 
32'd711: dataIn1 = 32'd13; 
32'd712: dataIn1 = 32'd24; 
32'd713: dataIn1 = 32'd23; 
32'd714: dataIn1 = 32'd24; 
32'd715: dataIn1 = 32'd14; 
32'd716: dataIn1 = 32'd28; 
32'd717: dataIn1 = 32'd31; 
32'd718: dataIn1 = 32'd19; 
32'd719: dataIn1 = 32'd10; 
32'd720: dataIn1 = 32'd19; 
32'd721: dataIn1 = 32'd15; 
32'd722: dataIn1 = 32'd18; 
32'd723: dataIn1 = 32'd24; 
32'd724: dataIn1 = 32'd31; 
32'd725: dataIn1 = 32'd13; 
32'd726: dataIn1 = 32'd30; 
32'd727: dataIn1 = 32'd24; 
32'd728: dataIn1 = 32'd16; 
32'd729: dataIn1 = 32'd21; 
32'd730: dataIn1 = 32'd8; 
32'd731: dataIn1 = 32'd24; 
32'd732: dataIn1 = 32'd11; 
32'd733: dataIn1 = 32'd28; 
32'd734: dataIn1 = 32'd19; 
32'd735: dataIn1 = 32'd10; 
32'd736: dataIn1 = 32'd24; 
32'd737: dataIn1 = 32'd13; 
32'd738: dataIn1 = 32'd25; 
32'd739: dataIn1 = 32'd21; 
32'd740: dataIn1 = 32'd2; 
32'd741: dataIn1 = 32'd9; 
32'd742: dataIn1 = 32'd9; 
32'd743: dataIn1 = 32'd9; 
32'd744: dataIn1 = 32'd22; 
32'd745: dataIn1 = 32'd0; 
32'd746: dataIn1 = 32'd23; 
32'd747: dataIn1 = 32'd26; 
32'd748: dataIn1 = 32'd23; 
32'd749: dataIn1 = 32'd28; 
32'd750: dataIn1 = 32'd7; 
32'd751: dataIn1 = 32'd11; 
32'd752: dataIn1 = 32'd31; 
32'd753: dataIn1 = 32'd25; 
32'd754: dataIn1 = 32'd22; 
32'd755: dataIn1 = 32'd23; 
32'd756: dataIn1 = 32'd24; 
32'd757: dataIn1 = 32'd14; 
32'd758: dataIn1 = 32'd3; 
32'd759: dataIn1 = 32'd14; 
32'd760: dataIn1 = 32'd9; 
32'd761: dataIn1 = 32'd21; 
32'd762: dataIn1 = 32'd23; 
32'd763: dataIn1 = 32'd0; 
32'd764: dataIn1 = 32'd4; 
32'd765: dataIn1 = 32'd27; 
32'd766: dataIn1 = 32'd22; 
32'd767: dataIn1 = 32'd8; 
32'd768: dataIn1 = 32'd7; 
32'd769: dataIn1 = 32'd13; 
32'd770: dataIn1 = 32'd8; 
32'd771: dataIn1 = 32'd30; 
32'd772: dataIn1 = 32'd3; 
32'd773: dataIn1 = 32'd30; 
32'd774: dataIn1 = 32'd11; 
32'd775: dataIn1 = 32'd15; 
32'd776: dataIn1 = 32'd31; 
32'd777: dataIn1 = 32'd25; 
32'd778: dataIn1 = 32'd22; 
32'd779: dataIn1 = 32'd25; 
32'd780: dataIn1 = 32'd13; 
32'd781: dataIn1 = 32'd21; 
32'd782: dataIn1 = 32'd12; 
32'd783: dataIn1 = 32'd29; 
32'd784: dataIn1 = 32'd15; 
32'd785: dataIn1 = 32'd12; 
32'd786: dataIn1 = 32'd11; 
32'd787: dataIn1 = 32'd5; 
32'd788: dataIn1 = 32'd7; 
32'd789: dataIn1 = 32'd23; 
32'd790: dataIn1 = 32'd18; 
32'd791: dataIn1 = 32'd2; 
32'd792: dataIn1 = 32'd10; 
32'd793: dataIn1 = 32'd26; 
32'd794: dataIn1 = 32'd20; 
32'd795: dataIn1 = 32'd16; 
32'd796: dataIn1 = 32'd24; 
32'd797: dataIn1 = 32'd6; 
32'd798: dataIn1 = 32'd11; 
32'd799: dataIn1 = 32'd24; 
32'd800: dataIn1 = 32'd9; 
32'd801: dataIn1 = 32'd2; 
32'd802: dataIn1 = 32'd28; 
32'd803: dataIn1 = 32'd27; 
32'd804: dataIn1 = 32'd5; 
32'd805: dataIn1 = 32'd5; 
32'd806: dataIn1 = 32'd19; 
32'd807: dataIn1 = 32'd1; 
32'd808: dataIn1 = 32'd10; 
32'd809: dataIn1 = 32'd23; 
32'd810: dataIn1 = 32'd27; 
32'd811: dataIn1 = 32'd13; 
32'd812: dataIn1 = 32'd21; 
32'd813: dataIn1 = 32'd26; 
32'd814: dataIn1 = 32'd31; 
32'd815: dataIn1 = 32'd4; 
32'd816: dataIn1 = 32'd20; 
32'd817: dataIn1 = 32'd21; 
32'd818: dataIn1 = 32'd7; 
32'd819: dataIn1 = 32'd12; 
32'd820: dataIn1 = 32'd17; 
32'd821: dataIn1 = 32'd12; 
32'd822: dataIn1 = 32'd23; 
32'd823: dataIn1 = 32'd22; 
32'd824: dataIn1 = 32'd21; 
32'd825: dataIn1 = 32'd23; 
32'd826: dataIn1 = 32'd5; 
32'd827: dataIn1 = 32'd11; 
32'd828: dataIn1 = 32'd26; 
32'd829: dataIn1 = 32'd28; 
32'd830: dataIn1 = 32'd28; 
32'd831: dataIn1 = 32'd14; 
32'd832: dataIn1 = 32'd14; 
32'd833: dataIn1 = 32'd26; 
32'd834: dataIn1 = 32'd0; 
32'd835: dataIn1 = 32'd18; 
32'd836: dataIn1 = 32'd21; 
32'd837: dataIn1 = 32'd8; 
32'd838: dataIn1 = 32'd26; 
32'd839: dataIn1 = 32'd5; 
32'd840: dataIn1 = 32'd0; 
32'd841: dataIn1 = 32'd20; 
32'd842: dataIn1 = 32'd11; 
32'd843: dataIn1 = 32'd28; 
32'd844: dataIn1 = 32'd26; 
32'd845: dataIn1 = 32'd1; 
32'd846: dataIn1 = 32'd22; 
32'd847: dataIn1 = 32'd6; 
32'd848: dataIn1 = 32'd22; 
32'd849: dataIn1 = 32'd31; 
32'd850: dataIn1 = 32'd16; 
32'd851: dataIn1 = 32'd17; 
32'd852: dataIn1 = 32'd15; 
32'd853: dataIn1 = 32'd31; 
32'd854: dataIn1 = 32'd31; 
32'd855: dataIn1 = 32'd20; 
32'd856: dataIn1 = 32'd16; 
32'd857: dataIn1 = 32'd7; 
32'd858: dataIn1 = 32'd2; 
32'd859: dataIn1 = 32'd26; 
32'd860: dataIn1 = 32'd19; 
32'd861: dataIn1 = 32'd25; 
32'd862: dataIn1 = 32'd23; 
32'd863: dataIn1 = 32'd4; 
32'd864: dataIn1 = 32'd2; 
32'd865: dataIn1 = 32'd29; 
32'd866: dataIn1 = 32'd27; 
32'd867: dataIn1 = 32'd9; 
32'd868: dataIn1 = 32'd29; 
32'd869: dataIn1 = 32'd16; 
32'd870: dataIn1 = 32'd5; 
32'd871: dataIn1 = 32'd8; 
32'd872: dataIn1 = 32'd18; 
32'd873: dataIn1 = 32'd17; 
32'd874: dataIn1 = 32'd18; 
32'd875: dataIn1 = 32'd8; 
32'd876: dataIn1 = 32'd2; 
32'd877: dataIn1 = 32'd28; 
32'd878: dataIn1 = 32'd22; 
32'd879: dataIn1 = 32'd22; 
32'd880: dataIn1 = 32'd13; 
32'd881: dataIn1 = 32'd31; 
32'd882: dataIn1 = 32'd7; 
32'd883: dataIn1 = 32'd21; 
32'd884: dataIn1 = 32'd6; 
32'd885: dataIn1 = 32'd16; 
32'd886: dataIn1 = 32'd8; 
32'd887: dataIn1 = 32'd20; 
32'd888: dataIn1 = 32'd25; 
32'd889: dataIn1 = 32'd25; 
32'd890: dataIn1 = 32'd8; 
32'd891: dataIn1 = 32'd8; 
32'd892: dataIn1 = 32'd30; 
32'd893: dataIn1 = 32'd3; 
32'd894: dataIn1 = 32'd25; 
32'd895: dataIn1 = 32'd17; 
32'd896: dataIn1 = 32'd8; 
32'd897: dataIn1 = 32'd21; 
32'd898: dataIn1 = 32'd18; 
32'd899: dataIn1 = 32'd4; 
32'd900: dataIn1 = 32'd23; 
32'd901: dataIn1 = 32'd30; 
32'd902: dataIn1 = 32'd25; 
32'd903: dataIn1 = 32'd2; 
32'd904: dataIn1 = 32'd28; 
32'd905: dataIn1 = 32'd30; 
32'd906: dataIn1 = 32'd31; 
32'd907: dataIn1 = 32'd20; 
32'd908: dataIn1 = 32'd22; 
32'd909: dataIn1 = 32'd18; 
32'd910: dataIn1 = 32'd20; 
32'd911: dataIn1 = 32'd29; 
32'd912: dataIn1 = 32'd11; 
32'd913: dataIn1 = 32'd0; 
32'd914: dataIn1 = 32'd7; 
32'd915: dataIn1 = 32'd6; 
32'd916: dataIn1 = 32'd15; 
32'd917: dataIn1 = 32'd27; 
32'd918: dataIn1 = 32'd2; 
32'd919: dataIn1 = 32'd26; 
32'd920: dataIn1 = 32'd9; 
32'd921: dataIn1 = 32'd28; 
32'd922: dataIn1 = 32'd22; 
32'd923: dataIn1 = 32'd14; 
32'd924: dataIn1 = 32'd4; 
32'd925: dataIn1 = 32'd31; 
32'd926: dataIn1 = 32'd11; 
32'd927: dataIn1 = 32'd13; 
32'd928: dataIn1 = 32'd8; 
32'd929: dataIn1 = 32'd8; 
32'd930: dataIn1 = 32'd14; 
32'd931: dataIn1 = 32'd5; 
32'd932: dataIn1 = 32'd18; 
32'd933: dataIn1 = 32'd10; 
32'd934: dataIn1 = 32'd8; 
32'd935: dataIn1 = 32'd21; 
32'd936: dataIn1 = 32'd1; 
32'd937: dataIn1 = 32'd19; 
32'd938: dataIn1 = 32'd0; 
32'd939: dataIn1 = 32'd21; 
32'd940: dataIn1 = 32'd21; 
32'd941: dataIn1 = 32'd22; 
32'd942: dataIn1 = 32'd25; 
32'd943: dataIn1 = 32'd17; 
32'd944: dataIn1 = 32'd29; 
32'd945: dataIn1 = 32'd17; 
32'd946: dataIn1 = 32'd16; 
32'd947: dataIn1 = 32'd23; 
32'd948: dataIn1 = 32'd18; 
32'd949: dataIn1 = 32'd23; 
32'd950: dataIn1 = 32'd9; 
32'd951: dataIn1 = 32'd30; 
32'd952: dataIn1 = 32'd28; 
32'd953: dataIn1 = 32'd29; 
32'd954: dataIn1 = 32'd22; 
32'd955: dataIn1 = 32'd18; 
32'd956: dataIn1 = 32'd9; 
32'd957: dataIn1 = 32'd30; 
32'd958: dataIn1 = 32'd15; 
32'd959: dataIn1 = 32'd23; 
32'd960: dataIn1 = 32'd25; 
32'd961: dataIn1 = 32'd10; 
32'd962: dataIn1 = 32'd18; 
32'd963: dataIn1 = 32'd25; 
32'd964: dataIn1 = 32'd4; 
32'd965: dataIn1 = 32'd22; 
32'd966: dataIn1 = 32'd1; 
32'd967: dataIn1 = 32'd5; 
32'd968: dataIn1 = 32'd21; 
32'd969: dataIn1 = 32'd12; 
32'd970: dataIn1 = 32'd29; 
32'd971: dataIn1 = 32'd29; 
32'd972: dataIn1 = 32'd22; 
32'd973: dataIn1 = 32'd8; 
32'd974: dataIn1 = 32'd9; 
32'd975: dataIn1 = 32'd9; 
32'd976: dataIn1 = 32'd3; 
32'd977: dataIn1 = 32'd16; 
32'd978: dataIn1 = 32'd24; 
32'd979: dataIn1 = 32'd20; 
32'd980: dataIn1 = 32'd6; 
32'd981: dataIn1 = 32'd28; 
32'd982: dataIn1 = 32'd8; 
32'd983: dataIn1 = 32'd8; 
32'd984: dataIn1 = 32'd18; 
32'd985: dataIn1 = 32'd24; 
32'd986: dataIn1 = 32'd8; 
32'd987: dataIn1 = 32'd4; 
32'd988: dataIn1 = 32'd16; 
32'd989: dataIn1 = 32'd28; 
32'd990: dataIn1 = 32'd10; 
32'd991: dataIn1 = 32'd11; 
32'd992: dataIn1 = 32'd8; 
32'd993: dataIn1 = 32'd5; 
32'd994: dataIn1 = 32'd6; 
32'd995: dataIn1 = 32'd10; 
32'd996: dataIn1 = 32'd31; 
32'd997: dataIn1 = 32'd21; 
32'd998: dataIn1 = 32'd17; 
32'd999: dataIn1 = 32'd14; 
32'd1000: dataIn1 = 32'd27; 
32'd1001: dataIn1 = 32'd24; 
32'd1002: dataIn1 = 32'd8; 
32'd1003: dataIn1 = 32'd27; 
32'd1004: dataIn1 = 32'd9; 
32'd1005: dataIn1 = 32'd30; 
32'd1006: dataIn1 = 32'd16; 
32'd1007: dataIn1 = 32'd15; 
32'd1008: dataIn1 = 32'd21; 
32'd1009: dataIn1 = 32'd2; 
32'd1010: dataIn1 = 32'd7; 
32'd1011: dataIn1 = 32'd20; 
32'd1012: dataIn1 = 32'd14; 
32'd1013: dataIn1 = 32'd5; 
32'd1014: dataIn1 = 32'd8; 
32'd1015: dataIn1 = 32'd24; 
32'd1016: dataIn1 = 32'd17; 
32'd1017: dataIn1 = 32'd25; 
32'd1018: dataIn1 = 32'd10; 
32'd1019: dataIn1 = 32'd20; 
32'd1020: dataIn1 = 32'd19; 
32'd1021: dataIn1 = 32'd10; 
32'd1022: dataIn1 = 32'd10; 
32'd1023: dataIn1 = 32'd28; 
32'd1024: dataIn1 = 32'd11; 
32'd1025: dataIn1 = 32'd23; 
32'd1026: dataIn1 = 32'd8; 
32'd1027: dataIn1 = 32'd20; 
32'd1028: dataIn1 = 32'd15; 
32'd1029: dataIn1 = 32'd2; 
32'd1030: dataIn1 = 32'd6; 
32'd1031: dataIn1 = 32'd1; 
32'd1032: dataIn1 = 32'd12; 
32'd1033: dataIn1 = 32'd5; 
32'd1034: dataIn1 = 32'd31; 
32'd1035: dataIn1 = 32'd6; 
32'd1036: dataIn1 = 32'd0; 
32'd1037: dataIn1 = 32'd13; 
32'd1038: dataIn1 = 32'd9; 
32'd1039: dataIn1 = 32'd28; 
32'd1040: dataIn1 = 32'd17; 
32'd1041: dataIn1 = 32'd17; 
32'd1042: dataIn1 = 32'd6; 
32'd1043: dataIn1 = 32'd2; 
32'd1044: dataIn1 = 32'd16; 
32'd1045: dataIn1 = 32'd11; 
32'd1046: dataIn1 = 32'd15; 
32'd1047: dataIn1 = 32'd26; 
32'd1048: dataIn1 = 32'd8; 
32'd1049: dataIn1 = 32'd19; 
32'd1050: dataIn1 = 32'd1; 
32'd1051: dataIn1 = 32'd2; 
32'd1052: dataIn1 = 32'd22; 
32'd1053: dataIn1 = 32'd27; 
32'd1054: dataIn1 = 32'd25; 
32'd1055: dataIn1 = 32'd16; 
32'd1056: dataIn1 = 32'd25; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd9; 
32'd3: dataIn2 = 32'd60; 
32'd4: dataIn2 = 32'd13; 
32'd5: dataIn2 = 32'd23; 
32'd6: dataIn2 = 32'd86; 
32'd7: dataIn2 = 32'd11; 
32'd8: dataIn2 = 32'd67; 
32'd9: dataIn2 = 32'd95; 
32'd10: dataIn2 = 32'd2; 
32'd11: dataIn2 = 32'd84; 
32'd12: dataIn2 = 32'd6; 
32'd13: dataIn2 = 32'd94; 
32'd14: dataIn2 = 32'd49; 
32'd15: dataIn2 = 32'd95; 
32'd16: dataIn2 = 32'd17; 
32'd17: dataIn2 = 32'd97; 
32'd18: dataIn2 = 32'd49; 
32'd19: dataIn2 = 32'd64; 
32'd20: dataIn2 = 32'd39; 
32'd21: dataIn2 = 32'd1; 
32'd22: dataIn2 = 32'd19; 
32'd23: dataIn2 = 32'd41; 
32'd24: dataIn2 = 32'd22; 
32'd25: dataIn2 = 32'd69; 
32'd26: dataIn2 = 32'd42; 
32'd27: dataIn2 = 32'd80; 
32'd28: dataIn2 = 32'd26; 
32'd29: dataIn2 = 32'd46; 
32'd30: dataIn2 = 32'd86; 
32'd31: dataIn2 = 32'd12; 
32'd32: dataIn2 = 32'd30; 
32'd33: dataIn2 = 32'd3; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht_synth.vcd"); 
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
