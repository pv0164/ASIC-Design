//64x64 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 3686 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd330 ; 
  wdata_col_base = 32'd40160 ; 
  row_base = 32'd438460 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #384000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd438460: dataIn1 = 32'd0
; 
32'd438461: dataIn1 = 32'd58
; 
32'd438462: dataIn1 = 32'd112
; 
32'd438463: dataIn1 = 32'd166
; 
32'd438464: dataIn1 = 32'd218
; 
32'd438465: dataIn1 = 32'd270
; 
32'd438466: dataIn1 = 32'd324
; 
32'd438467: dataIn1 = 32'd383
; 
32'd438468: dataIn1 = 32'd435
; 
32'd438469: dataIn1 = 32'd492
; 
32'd438470: dataIn1 = 32'd545
; 
32'd438471: dataIn1 = 32'd596
; 
32'd438472: dataIn1 = 32'd652
; 
32'd438473: dataIn1 = 32'd707
; 
32'd438474: dataIn1 = 32'd763
; 
32'd438475: dataIn1 = 32'd816
; 
32'd438476: dataIn1 = 32'd865
; 
32'd438477: dataIn1 = 32'd921
; 
32'd438478: dataIn1 = 32'd977
; 
32'd438479: dataIn1 = 32'd1031
; 
32'd438480: dataIn1 = 32'd1084
; 
32'd438481: dataIn1 = 32'd1138
; 
32'd438482: dataIn1 = 32'd1195
; 
32'd438483: dataIn1 = 32'd1249
; 
32'd438484: dataIn1 = 32'd1300
; 
32'd438485: dataIn1 = 32'd1356
; 
32'd438486: dataIn1 = 32'd1410
; 
32'd438487: dataIn1 = 32'd1468
; 
32'd438488: dataIn1 = 32'd1522
; 
32'd438489: dataIn1 = 32'd1581
; 
32'd438490: dataIn1 = 32'd1634
; 
32'd438491: dataIn1 = 32'd1689
; 
32'd438492: dataIn1 = 32'd1738
; 
32'd438493: dataIn1 = 32'd1793
; 
32'd438494: dataIn1 = 32'd1843
; 
32'd438495: dataIn1 = 32'd1898
; 
32'd438496: dataIn1 = 32'd1954
; 
32'd438497: dataIn1 = 32'd2012
; 
32'd438498: dataIn1 = 32'd2067
; 
32'd438499: dataIn1 = 32'd2116
; 
32'd438500: dataIn1 = 32'd2173
; 
32'd438501: dataIn1 = 32'd2230
; 
32'd438502: dataIn1 = 32'd2290
; 
32'd438503: dataIn1 = 32'd2345
; 
32'd438504: dataIn1 = 32'd2400
; 
32'd438505: dataIn1 = 32'd2452
; 
32'd438506: dataIn1 = 32'd2512
; 
32'd438507: dataIn1 = 32'd2569
; 
32'd438508: dataIn1 = 32'd2624
; 
32'd438509: dataIn1 = 32'd2678
; 
32'd438510: dataIn1 = 32'd2734
; 
32'd438511: dataIn1 = 32'd2790
; 
32'd438512: dataIn1 = 32'd2835
; 
32'd438513: dataIn1 = 32'd2891
; 
32'd438514: dataIn1 = 32'd2943
; 
32'd438515: dataIn1 = 32'd3001
; 
32'd438516: dataIn1 = 32'd3059
; 
32'd438517: dataIn1 = 32'd3109
; 
32'd438518: dataIn1 = 32'd3166
; 
32'd438519: dataIn1 = 32'd3222
; 
32'd438520: dataIn1 = 32'd3279
; 
32'd438521: dataIn1 = 32'd3338
; 
32'd438522: dataIn1 = 32'd3399
; 
32'd438523: dataIn1 = 32'd3451
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd40160: dataIn1 = 32'd0
; 
32'd40161: dataIn1 = 32'd58
; 
32'd40162: dataIn1 = 32'd112
; 
32'd40163: dataIn1 = 32'd166
; 
32'd40164: dataIn1 = 32'd218
; 
32'd40165: dataIn1 = 32'd270
; 
32'd40166: dataIn1 = 32'd324
; 
32'd40167: dataIn1 = 32'd383
; 
32'd40168: dataIn1 = 32'd435
; 
32'd40169: dataIn1 = 32'd492
; 
32'd40170: dataIn1 = 32'd545
; 
32'd40171: dataIn1 = 32'd596
; 
32'd40172: dataIn1 = 32'd652
; 
32'd40173: dataIn1 = 32'd707
; 
32'd40174: dataIn1 = 32'd763
; 
32'd40175: dataIn1 = 32'd816
; 
32'd40176: dataIn1 = 32'd865
; 
32'd40177: dataIn1 = 32'd921
; 
32'd40178: dataIn1 = 32'd977
; 
32'd40179: dataIn1 = 32'd1031
; 
32'd40180: dataIn1 = 32'd1084
; 
32'd40181: dataIn1 = 32'd1138
; 
32'd40182: dataIn1 = 32'd1195
; 
32'd40183: dataIn1 = 32'd1249
; 
32'd40184: dataIn1 = 32'd1300
; 
32'd40185: dataIn1 = 32'd1356
; 
32'd40186: dataIn1 = 32'd1410
; 
32'd40187: dataIn1 = 32'd1468
; 
32'd40188: dataIn1 = 32'd1522
; 
32'd40189: dataIn1 = 32'd1581
; 
32'd40190: dataIn1 = 32'd1634
; 
32'd40191: dataIn1 = 32'd1689
; 
32'd40192: dataIn1 = 32'd1738
; 
32'd40193: dataIn1 = 32'd1793
; 
32'd40194: dataIn1 = 32'd1843
; 
32'd40195: dataIn1 = 32'd1898
; 
32'd40196: dataIn1 = 32'd1954
; 
32'd40197: dataIn1 = 32'd2012
; 
32'd40198: dataIn1 = 32'd2067
; 
32'd40199: dataIn1 = 32'd2116
; 
32'd40200: dataIn1 = 32'd2173
; 
32'd40201: dataIn1 = 32'd2230
; 
32'd40202: dataIn1 = 32'd2290
; 
32'd40203: dataIn1 = 32'd2345
; 
32'd40204: dataIn1 = 32'd2400
; 
32'd40205: dataIn1 = 32'd2452
; 
32'd40206: dataIn1 = 32'd2512
; 
32'd40207: dataIn1 = 32'd2569
; 
32'd40208: dataIn1 = 32'd2624
; 
32'd40209: dataIn1 = 32'd2678
; 
32'd40210: dataIn1 = 32'd2734
; 
32'd40211: dataIn1 = 32'd2790
; 
32'd40212: dataIn1 = 32'd2835
; 
32'd40213: dataIn1 = 32'd2891
; 
32'd40214: dataIn1 = 32'd2943
; 
32'd40215: dataIn1 = 32'd3001
; 
32'd40216: dataIn1 = 32'd3059
; 
32'd40217: dataIn1 = 32'd3109
; 
32'd40218: dataIn1 = 32'd3166
; 
32'd40219: dataIn1 = 32'd3222
; 
32'd40220: dataIn1 = 32'd3279
; 
32'd40221: dataIn1 = 32'd3338
; 
32'd40222: dataIn1 = 32'd3399
; 
32'd40223: dataIn1 = 32'd3451
; 
32'd40224: dataIn1 = 32'd3506
; 
32'd40225: dataIn1 = 32'd0
; 
32'd40226: dataIn1 = 32'd1
; 
32'd40227: dataIn1 = 32'd2
; 
32'd40228: dataIn1 = 32'd3
; 
32'd40229: dataIn1 = 32'd5
; 
32'd40230: dataIn1 = 32'd6
; 
32'd40231: dataIn1 = 32'd7
; 
32'd40232: dataIn1 = 32'd8
; 
32'd40233: dataIn1 = 32'd9
; 
32'd40234: dataIn1 = 32'd10
; 
32'd40235: dataIn1 = 32'd11
; 
32'd40236: dataIn1 = 32'd12
; 
32'd40237: dataIn1 = 32'd13
; 
32'd40238: dataIn1 = 32'd14
; 
32'd40239: dataIn1 = 32'd15
; 
32'd40240: dataIn1 = 32'd16
; 
32'd40241: dataIn1 = 32'd17
; 
32'd40242: dataIn1 = 32'd18
; 
32'd40243: dataIn1 = 32'd20
; 
32'd40244: dataIn1 = 32'd21
; 
32'd40245: dataIn1 = 32'd22
; 
32'd40246: dataIn1 = 32'd23
; 
32'd40247: dataIn1 = 32'd24
; 
32'd40248: dataIn1 = 32'd25
; 
32'd40249: dataIn1 = 32'd27
; 
32'd40250: dataIn1 = 32'd28
; 
32'd40251: dataIn1 = 32'd29
; 
32'd40252: dataIn1 = 32'd30
; 
32'd40253: dataIn1 = 32'd31
; 
32'd40254: dataIn1 = 32'd32
; 
32'd40255: dataIn1 = 32'd33
; 
32'd40256: dataIn1 = 32'd34
; 
32'd40257: dataIn1 = 32'd35
; 
32'd40258: dataIn1 = 32'd36
; 
32'd40259: dataIn1 = 32'd37
; 
32'd40260: dataIn1 = 32'd38
; 
32'd40261: dataIn1 = 32'd39
; 
32'd40262: dataIn1 = 32'd40
; 
32'd40263: dataIn1 = 32'd41
; 
32'd40264: dataIn1 = 32'd44
; 
32'd40265: dataIn1 = 32'd45
; 
32'd40266: dataIn1 = 32'd46
; 
32'd40267: dataIn1 = 32'd47
; 
32'd40268: dataIn1 = 32'd48
; 
32'd40269: dataIn1 = 32'd49
; 
32'd40270: dataIn1 = 32'd50
; 
32'd40271: dataIn1 = 32'd51
; 
32'd40272: dataIn1 = 32'd52
; 
32'd40273: dataIn1 = 32'd53
; 
32'd40274: dataIn1 = 32'd54
; 
32'd40275: dataIn1 = 32'd56
; 
32'd40276: dataIn1 = 32'd57
; 
32'd40277: dataIn1 = 32'd58
; 
32'd40278: dataIn1 = 32'd59
; 
32'd40279: dataIn1 = 32'd60
; 
32'd40280: dataIn1 = 32'd61
; 
32'd40281: dataIn1 = 32'd62
; 
32'd40282: dataIn1 = 32'd63
; 
32'd40283: dataIn1 = 32'd0
; 
32'd40284: dataIn1 = 32'd1
; 
32'd40285: dataIn1 = 32'd2
; 
32'd40286: dataIn1 = 32'd3
; 
32'd40287: dataIn1 = 32'd4
; 
32'd40288: dataIn1 = 32'd5
; 
32'd40289: dataIn1 = 32'd6
; 
32'd40290: dataIn1 = 32'd7
; 
32'd40291: dataIn1 = 32'd8
; 
32'd40292: dataIn1 = 32'd10
; 
32'd40293: dataIn1 = 32'd11
; 
32'd40294: dataIn1 = 32'd12
; 
32'd40295: dataIn1 = 32'd13
; 
32'd40296: dataIn1 = 32'd14
; 
32'd40297: dataIn1 = 32'd15
; 
32'd40298: dataIn1 = 32'd16
; 
32'd40299: dataIn1 = 32'd18
; 
32'd40300: dataIn1 = 32'd19
; 
32'd40301: dataIn1 = 32'd20
; 
32'd40302: dataIn1 = 32'd21
; 
32'd40303: dataIn1 = 32'd22
; 
32'd40304: dataIn1 = 32'd23
; 
32'd40305: dataIn1 = 32'd24
; 
32'd40306: dataIn1 = 32'd25
; 
32'd40307: dataIn1 = 32'd26
; 
32'd40308: dataIn1 = 32'd27
; 
32'd40309: dataIn1 = 32'd28
; 
32'd40310: dataIn1 = 32'd29
; 
32'd40311: dataIn1 = 32'd30
; 
32'd40312: dataIn1 = 32'd32
; 
32'd40313: dataIn1 = 32'd33
; 
32'd40314: dataIn1 = 32'd34
; 
32'd40315: dataIn1 = 32'd35
; 
32'd40316: dataIn1 = 32'd36
; 
32'd40317: dataIn1 = 32'd37
; 
32'd40318: dataIn1 = 32'd38
; 
32'd40319: dataIn1 = 32'd39
; 
32'd40320: dataIn1 = 32'd40
; 
32'd40321: dataIn1 = 32'd41
; 
32'd40322: dataIn1 = 32'd42
; 
32'd40323: dataIn1 = 32'd45
; 
32'd40324: dataIn1 = 32'd46
; 
32'd40325: dataIn1 = 32'd47
; 
32'd40326: dataIn1 = 32'd48
; 
32'd40327: dataIn1 = 32'd50
; 
32'd40328: dataIn1 = 32'd51
; 
32'd40329: dataIn1 = 32'd52
; 
32'd40330: dataIn1 = 32'd53
; 
32'd40331: dataIn1 = 32'd54
; 
32'd40332: dataIn1 = 32'd55
; 
32'd40333: dataIn1 = 32'd57
; 
32'd40334: dataIn1 = 32'd58
; 
32'd40335: dataIn1 = 32'd60
; 
32'd40336: dataIn1 = 32'd63
; 
32'd40337: dataIn1 = 32'd1
; 
32'd40338: dataIn1 = 32'd2
; 
32'd40339: dataIn1 = 32'd3
; 
32'd40340: dataIn1 = 32'd4
; 
32'd40341: dataIn1 = 32'd5
; 
32'd40342: dataIn1 = 32'd7
; 
32'd40343: dataIn1 = 32'd9
; 
32'd40344: dataIn1 = 32'd10
; 
32'd40345: dataIn1 = 32'd12
; 
32'd40346: dataIn1 = 32'd14
; 
32'd40347: dataIn1 = 32'd15
; 
32'd40348: dataIn1 = 32'd16
; 
32'd40349: dataIn1 = 32'd17
; 
32'd40350: dataIn1 = 32'd18
; 
32'd40351: dataIn1 = 32'd19
; 
32'd40352: dataIn1 = 32'd20
; 
32'd40353: dataIn1 = 32'd23
; 
32'd40354: dataIn1 = 32'd24
; 
32'd40355: dataIn1 = 32'd25
; 
32'd40356: dataIn1 = 32'd26
; 
32'd40357: dataIn1 = 32'd27
; 
32'd40358: dataIn1 = 32'd28
; 
32'd40359: dataIn1 = 32'd29
; 
32'd40360: dataIn1 = 32'd30
; 
32'd40361: dataIn1 = 32'd31
; 
32'd40362: dataIn1 = 32'd32
; 
32'd40363: dataIn1 = 32'd33
; 
32'd40364: dataIn1 = 32'd34
; 
32'd40365: dataIn1 = 32'd35
; 
32'd40366: dataIn1 = 32'd36
; 
32'd40367: dataIn1 = 32'd38
; 
32'd40368: dataIn1 = 32'd39
; 
32'd40369: dataIn1 = 32'd41
; 
32'd40370: dataIn1 = 32'd42
; 
32'd40371: dataIn1 = 32'd43
; 
32'd40372: dataIn1 = 32'd44
; 
32'd40373: dataIn1 = 32'd45
; 
32'd40374: dataIn1 = 32'd46
; 
32'd40375: dataIn1 = 32'd47
; 
32'd40376: dataIn1 = 32'd48
; 
32'd40377: dataIn1 = 32'd49
; 
32'd40378: dataIn1 = 32'd50
; 
32'd40379: dataIn1 = 32'd51
; 
32'd40380: dataIn1 = 32'd52
; 
32'd40381: dataIn1 = 32'd53
; 
32'd40382: dataIn1 = 32'd54
; 
32'd40383: dataIn1 = 32'd55
; 
32'd40384: dataIn1 = 32'd56
; 
32'd40385: dataIn1 = 32'd58
; 
32'd40386: dataIn1 = 32'd59
; 
32'd40387: dataIn1 = 32'd60
; 
32'd40388: dataIn1 = 32'd61
; 
32'd40389: dataIn1 = 32'd62
; 
32'd40390: dataIn1 = 32'd63
; 
32'd40391: dataIn1 = 32'd0
; 
32'd40392: dataIn1 = 32'd1
; 
32'd40393: dataIn1 = 32'd3
; 
32'd40394: dataIn1 = 32'd5
; 
32'd40395: dataIn1 = 32'd6
; 
32'd40396: dataIn1 = 32'd7
; 
32'd40397: dataIn1 = 32'd8
; 
32'd40398: dataIn1 = 32'd9
; 
32'd40399: dataIn1 = 32'd10
; 
32'd40400: dataIn1 = 32'd11
; 
32'd40401: dataIn1 = 32'd12
; 
32'd40402: dataIn1 = 32'd13
; 
32'd40403: dataIn1 = 32'd14
; 
32'd40404: dataIn1 = 32'd15
; 
32'd40405: dataIn1 = 32'd16
; 
32'd40406: dataIn1 = 32'd17
; 
32'd40407: dataIn1 = 32'd18
; 
32'd40408: dataIn1 = 32'd19
; 
32'd40409: dataIn1 = 32'd20
; 
32'd40410: dataIn1 = 32'd21
; 
32'd40411: dataIn1 = 32'd22
; 
32'd40412: dataIn1 = 32'd23
; 
32'd40413: dataIn1 = 32'd24
; 
32'd40414: dataIn1 = 32'd26
; 
32'd40415: dataIn1 = 32'd27
; 
32'd40416: dataIn1 = 32'd28
; 
32'd40417: dataIn1 = 32'd30
; 
32'd40418: dataIn1 = 32'd31
; 
32'd40419: dataIn1 = 32'd32
; 
32'd40420: dataIn1 = 32'd33
; 
32'd40421: dataIn1 = 32'd34
; 
32'd40422: dataIn1 = 32'd35
; 
32'd40423: dataIn1 = 32'd36
; 
32'd40424: dataIn1 = 32'd37
; 
32'd40425: dataIn1 = 32'd39
; 
32'd40426: dataIn1 = 32'd40
; 
32'd40427: dataIn1 = 32'd41
; 
32'd40428: dataIn1 = 32'd42
; 
32'd40429: dataIn1 = 32'd43
; 
32'd40430: dataIn1 = 32'd44
; 
32'd40431: dataIn1 = 32'd45
; 
32'd40432: dataIn1 = 32'd47
; 
32'd40433: dataIn1 = 32'd50
; 
32'd40434: dataIn1 = 32'd51
; 
32'd40435: dataIn1 = 32'd52
; 
32'd40436: dataIn1 = 32'd53
; 
32'd40437: dataIn1 = 32'd54
; 
32'd40438: dataIn1 = 32'd55
; 
32'd40439: dataIn1 = 32'd56
; 
32'd40440: dataIn1 = 32'd59
; 
32'd40441: dataIn1 = 32'd61
; 
32'd40442: dataIn1 = 32'd62
; 
32'd40443: dataIn1 = 32'd0
; 
32'd40444: dataIn1 = 32'd2
; 
32'd40445: dataIn1 = 32'd3
; 
32'd40446: dataIn1 = 32'd4
; 
32'd40447: dataIn1 = 32'd5
; 
32'd40448: dataIn1 = 32'd6
; 
32'd40449: dataIn1 = 32'd8
; 
32'd40450: dataIn1 = 32'd9
; 
32'd40451: dataIn1 = 32'd10
; 
32'd40452: dataIn1 = 32'd12
; 
32'd40453: dataIn1 = 32'd13
; 
32'd40454: dataIn1 = 32'd14
; 
32'd40455: dataIn1 = 32'd15
; 
32'd40456: dataIn1 = 32'd16
; 
32'd40457: dataIn1 = 32'd17
; 
32'd40458: dataIn1 = 32'd18
; 
32'd40459: dataIn1 = 32'd20
; 
32'd40460: dataIn1 = 32'd21
; 
32'd40461: dataIn1 = 32'd23
; 
32'd40462: dataIn1 = 32'd25
; 
32'd40463: dataIn1 = 32'd27
; 
32'd40464: dataIn1 = 32'd28
; 
32'd40465: dataIn1 = 32'd29
; 
32'd40466: dataIn1 = 32'd30
; 
32'd40467: dataIn1 = 32'd31
; 
32'd40468: dataIn1 = 32'd32
; 
32'd40469: dataIn1 = 32'd33
; 
32'd40470: dataIn1 = 32'd34
; 
32'd40471: dataIn1 = 32'd35
; 
32'd40472: dataIn1 = 32'd37
; 
32'd40473: dataIn1 = 32'd38
; 
32'd40474: dataIn1 = 32'd39
; 
32'd40475: dataIn1 = 32'd40
; 
32'd40476: dataIn1 = 32'd41
; 
32'd40477: dataIn1 = 32'd42
; 
32'd40478: dataIn1 = 32'd43
; 
32'd40479: dataIn1 = 32'd44
; 
32'd40480: dataIn1 = 32'd45
; 
32'd40481: dataIn1 = 32'd48
; 
32'd40482: dataIn1 = 32'd49
; 
32'd40483: dataIn1 = 32'd50
; 
32'd40484: dataIn1 = 32'd51
; 
32'd40485: dataIn1 = 32'd52
; 
32'd40486: dataIn1 = 32'd54
; 
32'd40487: dataIn1 = 32'd55
; 
32'd40488: dataIn1 = 32'd56
; 
32'd40489: dataIn1 = 32'd57
; 
32'd40490: dataIn1 = 32'd58
; 
32'd40491: dataIn1 = 32'd59
; 
32'd40492: dataIn1 = 32'd60
; 
32'd40493: dataIn1 = 32'd62
; 
32'd40494: dataIn1 = 32'd63
; 
32'd40495: dataIn1 = 32'd0
; 
32'd40496: dataIn1 = 32'd1
; 
32'd40497: dataIn1 = 32'd2
; 
32'd40498: dataIn1 = 32'd3
; 
32'd40499: dataIn1 = 32'd4
; 
32'd40500: dataIn1 = 32'd5
; 
32'd40501: dataIn1 = 32'd7
; 
32'd40502: dataIn1 = 32'd9
; 
32'd40503: dataIn1 = 32'd10
; 
32'd40504: dataIn1 = 32'd11
; 
32'd40505: dataIn1 = 32'd12
; 
32'd40506: dataIn1 = 32'd13
; 
32'd40507: dataIn1 = 32'd15
; 
32'd40508: dataIn1 = 32'd16
; 
32'd40509: dataIn1 = 32'd18
; 
32'd40510: dataIn1 = 32'd19
; 
32'd40511: dataIn1 = 32'd20
; 
32'd40512: dataIn1 = 32'd21
; 
32'd40513: dataIn1 = 32'd23
; 
32'd40514: dataIn1 = 32'd24
; 
32'd40515: dataIn1 = 32'd25
; 
32'd40516: dataIn1 = 32'd26
; 
32'd40517: dataIn1 = 32'd27
; 
32'd40518: dataIn1 = 32'd28
; 
32'd40519: dataIn1 = 32'd29
; 
32'd40520: dataIn1 = 32'd30
; 
32'd40521: dataIn1 = 32'd31
; 
32'd40522: dataIn1 = 32'd32
; 
32'd40523: dataIn1 = 32'd33
; 
32'd40524: dataIn1 = 32'd34
; 
32'd40525: dataIn1 = 32'd35
; 
32'd40526: dataIn1 = 32'd36
; 
32'd40527: dataIn1 = 32'd37
; 
32'd40528: dataIn1 = 32'd38
; 
32'd40529: dataIn1 = 32'd39
; 
32'd40530: dataIn1 = 32'd40
; 
32'd40531: dataIn1 = 32'd41
; 
32'd40532: dataIn1 = 32'd42
; 
32'd40533: dataIn1 = 32'd43
; 
32'd40534: dataIn1 = 32'd45
; 
32'd40535: dataIn1 = 32'd46
; 
32'd40536: dataIn1 = 32'd47
; 
32'd40537: dataIn1 = 32'd48
; 
32'd40538: dataIn1 = 32'd49
; 
32'd40539: dataIn1 = 32'd51
; 
32'd40540: dataIn1 = 32'd54
; 
32'd40541: dataIn1 = 32'd55
; 
32'd40542: dataIn1 = 32'd56
; 
32'd40543: dataIn1 = 32'd58
; 
32'd40544: dataIn1 = 32'd59
; 
32'd40545: dataIn1 = 32'd60
; 
32'd40546: dataIn1 = 32'd61
; 
32'd40547: dataIn1 = 32'd62
; 
32'd40548: dataIn1 = 32'd63
; 
32'd40549: dataIn1 = 32'd1
; 
32'd40550: dataIn1 = 32'd2
; 
32'd40551: dataIn1 = 32'd3
; 
32'd40552: dataIn1 = 32'd4
; 
32'd40553: dataIn1 = 32'd5
; 
32'd40554: dataIn1 = 32'd6
; 
32'd40555: dataIn1 = 32'd7
; 
32'd40556: dataIn1 = 32'd8
; 
32'd40557: dataIn1 = 32'd9
; 
32'd40558: dataIn1 = 32'd10
; 
32'd40559: dataIn1 = 32'd11
; 
32'd40560: dataIn1 = 32'd12
; 
32'd40561: dataIn1 = 32'd13
; 
32'd40562: dataIn1 = 32'd14
; 
32'd40563: dataIn1 = 32'd15
; 
32'd40564: dataIn1 = 32'd16
; 
32'd40565: dataIn1 = 32'd17
; 
32'd40566: dataIn1 = 32'd18
; 
32'd40567: dataIn1 = 32'd19
; 
32'd40568: dataIn1 = 32'd20
; 
32'd40569: dataIn1 = 32'd21
; 
32'd40570: dataIn1 = 32'd22
; 
32'd40571: dataIn1 = 32'd23
; 
32'd40572: dataIn1 = 32'd24
; 
32'd40573: dataIn1 = 32'd25
; 
32'd40574: dataIn1 = 32'd26
; 
32'd40575: dataIn1 = 32'd27
; 
32'd40576: dataIn1 = 32'd28
; 
32'd40577: dataIn1 = 32'd30
; 
32'd40578: dataIn1 = 32'd31
; 
32'd40579: dataIn1 = 32'd32
; 
32'd40580: dataIn1 = 32'd33
; 
32'd40581: dataIn1 = 32'd34
; 
32'd40582: dataIn1 = 32'd35
; 
32'd40583: dataIn1 = 32'd36
; 
32'd40584: dataIn1 = 32'd37
; 
32'd40585: dataIn1 = 32'd38
; 
32'd40586: dataIn1 = 32'd39
; 
32'd40587: dataIn1 = 32'd40
; 
32'd40588: dataIn1 = 32'd41
; 
32'd40589: dataIn1 = 32'd43
; 
32'd40590: dataIn1 = 32'd44
; 
32'd40591: dataIn1 = 32'd45
; 
32'd40592: dataIn1 = 32'd46
; 
32'd40593: dataIn1 = 32'd47
; 
32'd40594: dataIn1 = 32'd48
; 
32'd40595: dataIn1 = 32'd50
; 
32'd40596: dataIn1 = 32'd51
; 
32'd40597: dataIn1 = 32'd52
; 
32'd40598: dataIn1 = 32'd53
; 
32'd40599: dataIn1 = 32'd54
; 
32'd40600: dataIn1 = 32'd55
; 
32'd40601: dataIn1 = 32'd56
; 
32'd40602: dataIn1 = 32'd57
; 
32'd40603: dataIn1 = 32'd58
; 
32'd40604: dataIn1 = 32'd59
; 
32'd40605: dataIn1 = 32'd60
; 
32'd40606: dataIn1 = 32'd61
; 
32'd40607: dataIn1 = 32'd63
; 
32'd40608: dataIn1 = 32'd0
; 
32'd40609: dataIn1 = 32'd3
; 
32'd40610: dataIn1 = 32'd4
; 
32'd40611: dataIn1 = 32'd5
; 
32'd40612: dataIn1 = 32'd6
; 
32'd40613: dataIn1 = 32'd7
; 
32'd40614: dataIn1 = 32'd8
; 
32'd40615: dataIn1 = 32'd9
; 
32'd40616: dataIn1 = 32'd10
; 
32'd40617: dataIn1 = 32'd12
; 
32'd40618: dataIn1 = 32'd13
; 
32'd40619: dataIn1 = 32'd14
; 
32'd40620: dataIn1 = 32'd15
; 
32'd40621: dataIn1 = 32'd16
; 
32'd40622: dataIn1 = 32'd17
; 
32'd40623: dataIn1 = 32'd18
; 
32'd40624: dataIn1 = 32'd20
; 
32'd40625: dataIn1 = 32'd21
; 
32'd40626: dataIn1 = 32'd22
; 
32'd40627: dataIn1 = 32'd24
; 
32'd40628: dataIn1 = 32'd25
; 
32'd40629: dataIn1 = 32'd26
; 
32'd40630: dataIn1 = 32'd27
; 
32'd40631: dataIn1 = 32'd28
; 
32'd40632: dataIn1 = 32'd29
; 
32'd40633: dataIn1 = 32'd31
; 
32'd40634: dataIn1 = 32'd32
; 
32'd40635: dataIn1 = 32'd33
; 
32'd40636: dataIn1 = 32'd34
; 
32'd40637: dataIn1 = 32'd35
; 
32'd40638: dataIn1 = 32'd36
; 
32'd40639: dataIn1 = 32'd37
; 
32'd40640: dataIn1 = 32'd38
; 
32'd40641: dataIn1 = 32'd39
; 
32'd40642: dataIn1 = 32'd40
; 
32'd40643: dataIn1 = 32'd41
; 
32'd40644: dataIn1 = 32'd42
; 
32'd40645: dataIn1 = 32'd43
; 
32'd40646: dataIn1 = 32'd44
; 
32'd40647: dataIn1 = 32'd47
; 
32'd40648: dataIn1 = 32'd49
; 
32'd40649: dataIn1 = 32'd50
; 
32'd40650: dataIn1 = 32'd51
; 
32'd40651: dataIn1 = 32'd52
; 
32'd40652: dataIn1 = 32'd53
; 
32'd40653: dataIn1 = 32'd54
; 
32'd40654: dataIn1 = 32'd55
; 
32'd40655: dataIn1 = 32'd56
; 
32'd40656: dataIn1 = 32'd57
; 
32'd40657: dataIn1 = 32'd60
; 
32'd40658: dataIn1 = 32'd62
; 
32'd40659: dataIn1 = 32'd63
; 
32'd40660: dataIn1 = 32'd0
; 
32'd40661: dataIn1 = 32'd1
; 
32'd40662: dataIn1 = 32'd2
; 
32'd40663: dataIn1 = 32'd4
; 
32'd40664: dataIn1 = 32'd5
; 
32'd40665: dataIn1 = 32'd6
; 
32'd40666: dataIn1 = 32'd7
; 
32'd40667: dataIn1 = 32'd8
; 
32'd40668: dataIn1 = 32'd9
; 
32'd40669: dataIn1 = 32'd10
; 
32'd40670: dataIn1 = 32'd11
; 
32'd40671: dataIn1 = 32'd12
; 
32'd40672: dataIn1 = 32'd13
; 
32'd40673: dataIn1 = 32'd14
; 
32'd40674: dataIn1 = 32'd15
; 
32'd40675: dataIn1 = 32'd16
; 
32'd40676: dataIn1 = 32'd17
; 
32'd40677: dataIn1 = 32'd18
; 
32'd40678: dataIn1 = 32'd20
; 
32'd40679: dataIn1 = 32'd21
; 
32'd40680: dataIn1 = 32'd22
; 
32'd40681: dataIn1 = 32'd23
; 
32'd40682: dataIn1 = 32'd24
; 
32'd40683: dataIn1 = 32'd25
; 
32'd40684: dataIn1 = 32'd26
; 
32'd40685: dataIn1 = 32'd27
; 
32'd40686: dataIn1 = 32'd28
; 
32'd40687: dataIn1 = 32'd29
; 
32'd40688: dataIn1 = 32'd30
; 
32'd40689: dataIn1 = 32'd31
; 
32'd40690: dataIn1 = 32'd32
; 
32'd40691: dataIn1 = 32'd34
; 
32'd40692: dataIn1 = 32'd35
; 
32'd40693: dataIn1 = 32'd36
; 
32'd40694: dataIn1 = 32'd37
; 
32'd40695: dataIn1 = 32'd39
; 
32'd40696: dataIn1 = 32'd40
; 
32'd40697: dataIn1 = 32'd41
; 
32'd40698: dataIn1 = 32'd42
; 
32'd40699: dataIn1 = 32'd43
; 
32'd40700: dataIn1 = 32'd44
; 
32'd40701: dataIn1 = 32'd45
; 
32'd40702: dataIn1 = 32'd46
; 
32'd40703: dataIn1 = 32'd48
; 
32'd40704: dataIn1 = 32'd50
; 
32'd40705: dataIn1 = 32'd51
; 
32'd40706: dataIn1 = 32'd52
; 
32'd40707: dataIn1 = 32'd53
; 
32'd40708: dataIn1 = 32'd54
; 
32'd40709: dataIn1 = 32'd55
; 
32'd40710: dataIn1 = 32'd56
; 
32'd40711: dataIn1 = 32'd58
; 
32'd40712: dataIn1 = 32'd59
; 
32'd40713: dataIn1 = 32'd60
; 
32'd40714: dataIn1 = 32'd61
; 
32'd40715: dataIn1 = 32'd62
; 
32'd40716: dataIn1 = 32'd63
; 
32'd40717: dataIn1 = 32'd0
; 
32'd40718: dataIn1 = 32'd2
; 
32'd40719: dataIn1 = 32'd3
; 
32'd40720: dataIn1 = 32'd4
; 
32'd40721: dataIn1 = 32'd5
; 
32'd40722: dataIn1 = 32'd6
; 
32'd40723: dataIn1 = 32'd7
; 
32'd40724: dataIn1 = 32'd8
; 
32'd40725: dataIn1 = 32'd9
; 
32'd40726: dataIn1 = 32'd11
; 
32'd40727: dataIn1 = 32'd12
; 
32'd40728: dataIn1 = 32'd13
; 
32'd40729: dataIn1 = 32'd14
; 
32'd40730: dataIn1 = 32'd15
; 
32'd40731: dataIn1 = 32'd16
; 
32'd40732: dataIn1 = 32'd17
; 
32'd40733: dataIn1 = 32'd18
; 
32'd40734: dataIn1 = 32'd19
; 
32'd40735: dataIn1 = 32'd20
; 
32'd40736: dataIn1 = 32'd21
; 
32'd40737: dataIn1 = 32'd22
; 
32'd40738: dataIn1 = 32'd23
; 
32'd40739: dataIn1 = 32'd25
; 
32'd40740: dataIn1 = 32'd26
; 
32'd40741: dataIn1 = 32'd27
; 
32'd40742: dataIn1 = 32'd28
; 
32'd40743: dataIn1 = 32'd29
; 
32'd40744: dataIn1 = 32'd30
; 
32'd40745: dataIn1 = 32'd31
; 
32'd40746: dataIn1 = 32'd32
; 
32'd40747: dataIn1 = 32'd34
; 
32'd40748: dataIn1 = 32'd35
; 
32'd40749: dataIn1 = 32'd36
; 
32'd40750: dataIn1 = 32'd37
; 
32'd40751: dataIn1 = 32'd38
; 
32'd40752: dataIn1 = 32'd39
; 
32'd40753: dataIn1 = 32'd41
; 
32'd40754: dataIn1 = 32'd42
; 
32'd40755: dataIn1 = 32'd43
; 
32'd40756: dataIn1 = 32'd46
; 
32'd40757: dataIn1 = 32'd47
; 
32'd40758: dataIn1 = 32'd48
; 
32'd40759: dataIn1 = 32'd49
; 
32'd40760: dataIn1 = 32'd50
; 
32'd40761: dataIn1 = 32'd52
; 
32'd40762: dataIn1 = 32'd53
; 
32'd40763: dataIn1 = 32'd54
; 
32'd40764: dataIn1 = 32'd55
; 
32'd40765: dataIn1 = 32'd58
; 
32'd40766: dataIn1 = 32'd59
; 
32'd40767: dataIn1 = 32'd60
; 
32'd40768: dataIn1 = 32'd61
; 
32'd40769: dataIn1 = 32'd63
; 
32'd40770: dataIn1 = 32'd1
; 
32'd40771: dataIn1 = 32'd2
; 
32'd40772: dataIn1 = 32'd3
; 
32'd40773: dataIn1 = 32'd4
; 
32'd40774: dataIn1 = 32'd5
; 
32'd40775: dataIn1 = 32'd6
; 
32'd40776: dataIn1 = 32'd7
; 
32'd40777: dataIn1 = 32'd8
; 
32'd40778: dataIn1 = 32'd9
; 
32'd40779: dataIn1 = 32'd10
; 
32'd40780: dataIn1 = 32'd12
; 
32'd40781: dataIn1 = 32'd13
; 
32'd40782: dataIn1 = 32'd17
; 
32'd40783: dataIn1 = 32'd18
; 
32'd40784: dataIn1 = 32'd19
; 
32'd40785: dataIn1 = 32'd21
; 
32'd40786: dataIn1 = 32'd22
; 
32'd40787: dataIn1 = 32'd24
; 
32'd40788: dataIn1 = 32'd25
; 
32'd40789: dataIn1 = 32'd26
; 
32'd40790: dataIn1 = 32'd27
; 
32'd40791: dataIn1 = 32'd28
; 
32'd40792: dataIn1 = 32'd29
; 
32'd40793: dataIn1 = 32'd30
; 
32'd40794: dataIn1 = 32'd31
; 
32'd40795: dataIn1 = 32'd32
; 
32'd40796: dataIn1 = 32'd33
; 
32'd40797: dataIn1 = 32'd34
; 
32'd40798: dataIn1 = 32'd35
; 
32'd40799: dataIn1 = 32'd38
; 
32'd40800: dataIn1 = 32'd41
; 
32'd40801: dataIn1 = 32'd42
; 
32'd40802: dataIn1 = 32'd43
; 
32'd40803: dataIn1 = 32'd44
; 
32'd40804: dataIn1 = 32'd45
; 
32'd40805: dataIn1 = 32'd46
; 
32'd40806: dataIn1 = 32'd47
; 
32'd40807: dataIn1 = 32'd48
; 
32'd40808: dataIn1 = 32'd49
; 
32'd40809: dataIn1 = 32'd50
; 
32'd40810: dataIn1 = 32'd51
; 
32'd40811: dataIn1 = 32'd52
; 
32'd40812: dataIn1 = 32'd54
; 
32'd40813: dataIn1 = 32'd55
; 
32'd40814: dataIn1 = 32'd56
; 
32'd40815: dataIn1 = 32'd57
; 
32'd40816: dataIn1 = 32'd59
; 
32'd40817: dataIn1 = 32'd60
; 
32'd40818: dataIn1 = 32'd61
; 
32'd40819: dataIn1 = 32'd62
; 
32'd40820: dataIn1 = 32'd63
; 
32'd40821: dataIn1 = 32'd2
; 
32'd40822: dataIn1 = 32'd3
; 
32'd40823: dataIn1 = 32'd4
; 
32'd40824: dataIn1 = 32'd5
; 
32'd40825: dataIn1 = 32'd6
; 
32'd40826: dataIn1 = 32'd7
; 
32'd40827: dataIn1 = 32'd8
; 
32'd40828: dataIn1 = 32'd9
; 
32'd40829: dataIn1 = 32'd10
; 
32'd40830: dataIn1 = 32'd11
; 
32'd40831: dataIn1 = 32'd12
; 
32'd40832: dataIn1 = 32'd13
; 
32'd40833: dataIn1 = 32'd15
; 
32'd40834: dataIn1 = 32'd16
; 
32'd40835: dataIn1 = 32'd17
; 
32'd40836: dataIn1 = 32'd18
; 
32'd40837: dataIn1 = 32'd19
; 
32'd40838: dataIn1 = 32'd20
; 
32'd40839: dataIn1 = 32'd22
; 
32'd40840: dataIn1 = 32'd23
; 
32'd40841: dataIn1 = 32'd24
; 
32'd40842: dataIn1 = 32'd25
; 
32'd40843: dataIn1 = 32'd26
; 
32'd40844: dataIn1 = 32'd27
; 
32'd40845: dataIn1 = 32'd28
; 
32'd40846: dataIn1 = 32'd29
; 
32'd40847: dataIn1 = 32'd30
; 
32'd40848: dataIn1 = 32'd31
; 
32'd40849: dataIn1 = 32'd32
; 
32'd40850: dataIn1 = 32'd33
; 
32'd40851: dataIn1 = 32'd35
; 
32'd40852: dataIn1 = 32'd36
; 
32'd40853: dataIn1 = 32'd37
; 
32'd40854: dataIn1 = 32'd38
; 
32'd40855: dataIn1 = 32'd39
; 
32'd40856: dataIn1 = 32'd40
; 
32'd40857: dataIn1 = 32'd41
; 
32'd40858: dataIn1 = 32'd43
; 
32'd40859: dataIn1 = 32'd45
; 
32'd40860: dataIn1 = 32'd46
; 
32'd40861: dataIn1 = 32'd47
; 
32'd40862: dataIn1 = 32'd48
; 
32'd40863: dataIn1 = 32'd49
; 
32'd40864: dataIn1 = 32'd50
; 
32'd40865: dataIn1 = 32'd51
; 
32'd40866: dataIn1 = 32'd52
; 
32'd40867: dataIn1 = 32'd54
; 
32'd40868: dataIn1 = 32'd55
; 
32'd40869: dataIn1 = 32'd56
; 
32'd40870: dataIn1 = 32'd57
; 
32'd40871: dataIn1 = 32'd58
; 
32'd40872: dataIn1 = 32'd59
; 
32'd40873: dataIn1 = 32'd60
; 
32'd40874: dataIn1 = 32'd61
; 
32'd40875: dataIn1 = 32'd62
; 
32'd40876: dataIn1 = 32'd63
; 
32'd40877: dataIn1 = 32'd1
; 
32'd40878: dataIn1 = 32'd2
; 
32'd40879: dataIn1 = 32'd3
; 
32'd40880: dataIn1 = 32'd4
; 
32'd40881: dataIn1 = 32'd5
; 
32'd40882: dataIn1 = 32'd6
; 
32'd40883: dataIn1 = 32'd7
; 
32'd40884: dataIn1 = 32'd8
; 
32'd40885: dataIn1 = 32'd9
; 
32'd40886: dataIn1 = 32'd11
; 
32'd40887: dataIn1 = 32'd12
; 
32'd40888: dataIn1 = 32'd13
; 
32'd40889: dataIn1 = 32'd14
; 
32'd40890: dataIn1 = 32'd16
; 
32'd40891: dataIn1 = 32'd17
; 
32'd40892: dataIn1 = 32'd18
; 
32'd40893: dataIn1 = 32'd19
; 
32'd40894: dataIn1 = 32'd20
; 
32'd40895: dataIn1 = 32'd21
; 
32'd40896: dataIn1 = 32'd22
; 
32'd40897: dataIn1 = 32'd23
; 
32'd40898: dataIn1 = 32'd24
; 
32'd40899: dataIn1 = 32'd26
; 
32'd40900: dataIn1 = 32'd28
; 
32'd40901: dataIn1 = 32'd29
; 
32'd40902: dataIn1 = 32'd31
; 
32'd40903: dataIn1 = 32'd32
; 
32'd40904: dataIn1 = 32'd33
; 
32'd40905: dataIn1 = 32'd34
; 
32'd40906: dataIn1 = 32'd35
; 
32'd40907: dataIn1 = 32'd36
; 
32'd40908: dataIn1 = 32'd37
; 
32'd40909: dataIn1 = 32'd38
; 
32'd40910: dataIn1 = 32'd40
; 
32'd40911: dataIn1 = 32'd41
; 
32'd40912: dataIn1 = 32'd42
; 
32'd40913: dataIn1 = 32'd44
; 
32'd40914: dataIn1 = 32'd45
; 
32'd40915: dataIn1 = 32'd46
; 
32'd40916: dataIn1 = 32'd47
; 
32'd40917: dataIn1 = 32'd48
; 
32'd40918: dataIn1 = 32'd49
; 
32'd40919: dataIn1 = 32'd50
; 
32'd40920: dataIn1 = 32'd51
; 
32'd40921: dataIn1 = 32'd52
; 
32'd40922: dataIn1 = 32'd53
; 
32'd40923: dataIn1 = 32'd54
; 
32'd40924: dataIn1 = 32'd55
; 
32'd40925: dataIn1 = 32'd56
; 
32'd40926: dataIn1 = 32'd57
; 
32'd40927: dataIn1 = 32'd58
; 
32'd40928: dataIn1 = 32'd59
; 
32'd40929: dataIn1 = 32'd60
; 
32'd40930: dataIn1 = 32'd61
; 
32'd40931: dataIn1 = 32'd62
; 
32'd40932: dataIn1 = 32'd0
; 
32'd40933: dataIn1 = 32'd1
; 
32'd40934: dataIn1 = 32'd2
; 
32'd40935: dataIn1 = 32'd3
; 
32'd40936: dataIn1 = 32'd4
; 
32'd40937: dataIn1 = 32'd5
; 
32'd40938: dataIn1 = 32'd6
; 
32'd40939: dataIn1 = 32'd7
; 
32'd40940: dataIn1 = 32'd8
; 
32'd40941: dataIn1 = 32'd9
; 
32'd40942: dataIn1 = 32'd10
; 
32'd40943: dataIn1 = 32'd11
; 
32'd40944: dataIn1 = 32'd12
; 
32'd40945: dataIn1 = 32'd13
; 
32'd40946: dataIn1 = 32'd15
; 
32'd40947: dataIn1 = 32'd16
; 
32'd40948: dataIn1 = 32'd18
; 
32'd40949: dataIn1 = 32'd19
; 
32'd40950: dataIn1 = 32'd20
; 
32'd40951: dataIn1 = 32'd21
; 
32'd40952: dataIn1 = 32'd22
; 
32'd40953: dataIn1 = 32'd24
; 
32'd40954: dataIn1 = 32'd25
; 
32'd40955: dataIn1 = 32'd26
; 
32'd40956: dataIn1 = 32'd29
; 
32'd40957: dataIn1 = 32'd30
; 
32'd40958: dataIn1 = 32'd31
; 
32'd40959: dataIn1 = 32'd33
; 
32'd40960: dataIn1 = 32'd34
; 
32'd40961: dataIn1 = 32'd35
; 
32'd40962: dataIn1 = 32'd36
; 
32'd40963: dataIn1 = 32'd37
; 
32'd40964: dataIn1 = 32'd38
; 
32'd40965: dataIn1 = 32'd39
; 
32'd40966: dataIn1 = 32'd40
; 
32'd40967: dataIn1 = 32'd41
; 
32'd40968: dataIn1 = 32'd42
; 
32'd40969: dataIn1 = 32'd43
; 
32'd40970: dataIn1 = 32'd45
; 
32'd40971: dataIn1 = 32'd46
; 
32'd40972: dataIn1 = 32'd47
; 
32'd40973: dataIn1 = 32'd49
; 
32'd40974: dataIn1 = 32'd50
; 
32'd40975: dataIn1 = 32'd51
; 
32'd40976: dataIn1 = 32'd52
; 
32'd40977: dataIn1 = 32'd53
; 
32'd40978: dataIn1 = 32'd54
; 
32'd40979: dataIn1 = 32'd55
; 
32'd40980: dataIn1 = 32'd56
; 
32'd40981: dataIn1 = 32'd57
; 
32'd40982: dataIn1 = 32'd58
; 
32'd40983: dataIn1 = 32'd59
; 
32'd40984: dataIn1 = 32'd60
; 
32'd40985: dataIn1 = 32'd61
; 
32'd40986: dataIn1 = 32'd62
; 
32'd40987: dataIn1 = 32'd63
; 
32'd40988: dataIn1 = 32'd0
; 
32'd40989: dataIn1 = 32'd1
; 
32'd40990: dataIn1 = 32'd2
; 
32'd40991: dataIn1 = 32'd3
; 
32'd40992: dataIn1 = 32'd5
; 
32'd40993: dataIn1 = 32'd6
; 
32'd40994: dataIn1 = 32'd7
; 
32'd40995: dataIn1 = 32'd8
; 
32'd40996: dataIn1 = 32'd9
; 
32'd40997: dataIn1 = 32'd10
; 
32'd40998: dataIn1 = 32'd11
; 
32'd40999: dataIn1 = 32'd13
; 
32'd41000: dataIn1 = 32'd14
; 
32'd41001: dataIn1 = 32'd16
; 
32'd41002: dataIn1 = 32'd17
; 
32'd41003: dataIn1 = 32'd21
; 
32'd41004: dataIn1 = 32'd22
; 
32'd41005: dataIn1 = 32'd23
; 
32'd41006: dataIn1 = 32'd24
; 
32'd41007: dataIn1 = 32'd25
; 
32'd41008: dataIn1 = 32'd26
; 
32'd41009: dataIn1 = 32'd27
; 
32'd41010: dataIn1 = 32'd28
; 
32'd41011: dataIn1 = 32'd31
; 
32'd41012: dataIn1 = 32'd32
; 
32'd41013: dataIn1 = 32'd33
; 
32'd41014: dataIn1 = 32'd34
; 
32'd41015: dataIn1 = 32'd36
; 
32'd41016: dataIn1 = 32'd37
; 
32'd41017: dataIn1 = 32'd38
; 
32'd41018: dataIn1 = 32'd40
; 
32'd41019: dataIn1 = 32'd41
; 
32'd41020: dataIn1 = 32'd42
; 
32'd41021: dataIn1 = 32'd43
; 
32'd41022: dataIn1 = 32'd44
; 
32'd41023: dataIn1 = 32'd45
; 
32'd41024: dataIn1 = 32'd46
; 
32'd41025: dataIn1 = 32'd47
; 
32'd41026: dataIn1 = 32'd48
; 
32'd41027: dataIn1 = 32'd49
; 
32'd41028: dataIn1 = 32'd50
; 
32'd41029: dataIn1 = 32'd51
; 
32'd41030: dataIn1 = 32'd52
; 
32'd41031: dataIn1 = 32'd53
; 
32'd41032: dataIn1 = 32'd54
; 
32'd41033: dataIn1 = 32'd55
; 
32'd41034: dataIn1 = 32'd56
; 
32'd41035: dataIn1 = 32'd57
; 
32'd41036: dataIn1 = 32'd59
; 
32'd41037: dataIn1 = 32'd60
; 
32'd41038: dataIn1 = 32'd61
; 
32'd41039: dataIn1 = 32'd62
; 
32'd41040: dataIn1 = 32'd63
; 
32'd41041: dataIn1 = 32'd0
; 
32'd41042: dataIn1 = 32'd1
; 
32'd41043: dataIn1 = 32'd2
; 
32'd41044: dataIn1 = 32'd4
; 
32'd41045: dataIn1 = 32'd6
; 
32'd41046: dataIn1 = 32'd7
; 
32'd41047: dataIn1 = 32'd9
; 
32'd41048: dataIn1 = 32'd10
; 
32'd41049: dataIn1 = 32'd11
; 
32'd41050: dataIn1 = 32'd12
; 
32'd41051: dataIn1 = 32'd13
; 
32'd41052: dataIn1 = 32'd14
; 
32'd41053: dataIn1 = 32'd15
; 
32'd41054: dataIn1 = 32'd18
; 
32'd41055: dataIn1 = 32'd19
; 
32'd41056: dataIn1 = 32'd20
; 
32'd41057: dataIn1 = 32'd21
; 
32'd41058: dataIn1 = 32'd22
; 
32'd41059: dataIn1 = 32'd23
; 
32'd41060: dataIn1 = 32'd24
; 
32'd41061: dataIn1 = 32'd25
; 
32'd41062: dataIn1 = 32'd28
; 
32'd41063: dataIn1 = 32'd29
; 
32'd41064: dataIn1 = 32'd31
; 
32'd41065: dataIn1 = 32'd33
; 
32'd41066: dataIn1 = 32'd34
; 
32'd41067: dataIn1 = 32'd35
; 
32'd41068: dataIn1 = 32'd36
; 
32'd41069: dataIn1 = 32'd37
; 
32'd41070: dataIn1 = 32'd38
; 
32'd41071: dataIn1 = 32'd40
; 
32'd41072: dataIn1 = 32'd41
; 
32'd41073: dataIn1 = 32'd42
; 
32'd41074: dataIn1 = 32'd43
; 
32'd41075: dataIn1 = 32'd45
; 
32'd41076: dataIn1 = 32'd46
; 
32'd41077: dataIn1 = 32'd49
; 
32'd41078: dataIn1 = 32'd50
; 
32'd41079: dataIn1 = 32'd51
; 
32'd41080: dataIn1 = 32'd52
; 
32'd41081: dataIn1 = 32'd54
; 
32'd41082: dataIn1 = 32'd55
; 
32'd41083: dataIn1 = 32'd56
; 
32'd41084: dataIn1 = 32'd57
; 
32'd41085: dataIn1 = 32'd58
; 
32'd41086: dataIn1 = 32'd60
; 
32'd41087: dataIn1 = 32'd61
; 
32'd41088: dataIn1 = 32'd62
; 
32'd41089: dataIn1 = 32'd63
; 
32'd41090: dataIn1 = 32'd0
; 
32'd41091: dataIn1 = 32'd1
; 
32'd41092: dataIn1 = 32'd2
; 
32'd41093: dataIn1 = 32'd3
; 
32'd41094: dataIn1 = 32'd4
; 
32'd41095: dataIn1 = 32'd5
; 
32'd41096: dataIn1 = 32'd7
; 
32'd41097: dataIn1 = 32'd8
; 
32'd41098: dataIn1 = 32'd9
; 
32'd41099: dataIn1 = 32'd10
; 
32'd41100: dataIn1 = 32'd11
; 
32'd41101: dataIn1 = 32'd12
; 
32'd41102: dataIn1 = 32'd14
; 
32'd41103: dataIn1 = 32'd15
; 
32'd41104: dataIn1 = 32'd16
; 
32'd41105: dataIn1 = 32'd17
; 
32'd41106: dataIn1 = 32'd18
; 
32'd41107: dataIn1 = 32'd19
; 
32'd41108: dataIn1 = 32'd20
; 
32'd41109: dataIn1 = 32'd21
; 
32'd41110: dataIn1 = 32'd22
; 
32'd41111: dataIn1 = 32'd24
; 
32'd41112: dataIn1 = 32'd25
; 
32'd41113: dataIn1 = 32'd26
; 
32'd41114: dataIn1 = 32'd27
; 
32'd41115: dataIn1 = 32'd29
; 
32'd41116: dataIn1 = 32'd30
; 
32'd41117: dataIn1 = 32'd31
; 
32'd41118: dataIn1 = 32'd32
; 
32'd41119: dataIn1 = 32'd33
; 
32'd41120: dataIn1 = 32'd34
; 
32'd41121: dataIn1 = 32'd35
; 
32'd41122: dataIn1 = 32'd36
; 
32'd41123: dataIn1 = 32'd38
; 
32'd41124: dataIn1 = 32'd39
; 
32'd41125: dataIn1 = 32'd40
; 
32'd41126: dataIn1 = 32'd41
; 
32'd41127: dataIn1 = 32'd42
; 
32'd41128: dataIn1 = 32'd43
; 
32'd41129: dataIn1 = 32'd44
; 
32'd41130: dataIn1 = 32'd45
; 
32'd41131: dataIn1 = 32'd46
; 
32'd41132: dataIn1 = 32'd47
; 
32'd41133: dataIn1 = 32'd48
; 
32'd41134: dataIn1 = 32'd50
; 
32'd41135: dataIn1 = 32'd51
; 
32'd41136: dataIn1 = 32'd54
; 
32'd41137: dataIn1 = 32'd55
; 
32'd41138: dataIn1 = 32'd56
; 
32'd41139: dataIn1 = 32'd57
; 
32'd41140: dataIn1 = 32'd58
; 
32'd41141: dataIn1 = 32'd59
; 
32'd41142: dataIn1 = 32'd60
; 
32'd41143: dataIn1 = 32'd61
; 
32'd41144: dataIn1 = 32'd62
; 
32'd41145: dataIn1 = 32'd63
; 
32'd41146: dataIn1 = 32'd0
; 
32'd41147: dataIn1 = 32'd1
; 
32'd41148: dataIn1 = 32'd2
; 
32'd41149: dataIn1 = 32'd3
; 
32'd41150: dataIn1 = 32'd4
; 
32'd41151: dataIn1 = 32'd6
; 
32'd41152: dataIn1 = 32'd7
; 
32'd41153: dataIn1 = 32'd8
; 
32'd41154: dataIn1 = 32'd9
; 
32'd41155: dataIn1 = 32'd10
; 
32'd41156: dataIn1 = 32'd11
; 
32'd41157: dataIn1 = 32'd12
; 
32'd41158: dataIn1 = 32'd13
; 
32'd41159: dataIn1 = 32'd14
; 
32'd41160: dataIn1 = 32'd15
; 
32'd41161: dataIn1 = 32'd16
; 
32'd41162: dataIn1 = 32'd17
; 
32'd41163: dataIn1 = 32'd18
; 
32'd41164: dataIn1 = 32'd19
; 
32'd41165: dataIn1 = 32'd20
; 
32'd41166: dataIn1 = 32'd21
; 
32'd41167: dataIn1 = 32'd24
; 
32'd41168: dataIn1 = 32'd25
; 
32'd41169: dataIn1 = 32'd29
; 
32'd41170: dataIn1 = 32'd30
; 
32'd41171: dataIn1 = 32'd31
; 
32'd41172: dataIn1 = 32'd32
; 
32'd41173: dataIn1 = 32'd33
; 
32'd41174: dataIn1 = 32'd34
; 
32'd41175: dataIn1 = 32'd35
; 
32'd41176: dataIn1 = 32'd36
; 
32'd41177: dataIn1 = 32'd37
; 
32'd41178: dataIn1 = 32'd38
; 
32'd41179: dataIn1 = 32'd39
; 
32'd41180: dataIn1 = 32'd40
; 
32'd41181: dataIn1 = 32'd41
; 
32'd41182: dataIn1 = 32'd42
; 
32'd41183: dataIn1 = 32'd43
; 
32'd41184: dataIn1 = 32'd44
; 
32'd41185: dataIn1 = 32'd45
; 
32'd41186: dataIn1 = 32'd46
; 
32'd41187: dataIn1 = 32'd47
; 
32'd41188: dataIn1 = 32'd49
; 
32'd41189: dataIn1 = 32'd50
; 
32'd41190: dataIn1 = 32'd51
; 
32'd41191: dataIn1 = 32'd52
; 
32'd41192: dataIn1 = 32'd53
; 
32'd41193: dataIn1 = 32'd54
; 
32'd41194: dataIn1 = 32'd55
; 
32'd41195: dataIn1 = 32'd56
; 
32'd41196: dataIn1 = 32'd57
; 
32'd41197: dataIn1 = 32'd58
; 
32'd41198: dataIn1 = 32'd59
; 
32'd41199: dataIn1 = 32'd61
; 
32'd41200: dataIn1 = 32'd62
; 
32'd41201: dataIn1 = 32'd63
; 
32'd41202: dataIn1 = 32'd1
; 
32'd41203: dataIn1 = 32'd2
; 
32'd41204: dataIn1 = 32'd3
; 
32'd41205: dataIn1 = 32'd4
; 
32'd41206: dataIn1 = 32'd6
; 
32'd41207: dataIn1 = 32'd7
; 
32'd41208: dataIn1 = 32'd8
; 
32'd41209: dataIn1 = 32'd9
; 
32'd41210: dataIn1 = 32'd10
; 
32'd41211: dataIn1 = 32'd12
; 
32'd41212: dataIn1 = 32'd13
; 
32'd41213: dataIn1 = 32'd14
; 
32'd41214: dataIn1 = 32'd15
; 
32'd41215: dataIn1 = 32'd16
; 
32'd41216: dataIn1 = 32'd17
; 
32'd41217: dataIn1 = 32'd18
; 
32'd41218: dataIn1 = 32'd19
; 
32'd41219: dataIn1 = 32'd20
; 
32'd41220: dataIn1 = 32'd21
; 
32'd41221: dataIn1 = 32'd22
; 
32'd41222: dataIn1 = 32'd23
; 
32'd41223: dataIn1 = 32'd24
; 
32'd41224: dataIn1 = 32'd25
; 
32'd41225: dataIn1 = 32'd26
; 
32'd41226: dataIn1 = 32'd27
; 
32'd41227: dataIn1 = 32'd28
; 
32'd41228: dataIn1 = 32'd29
; 
32'd41229: dataIn1 = 32'd30
; 
32'd41230: dataIn1 = 32'd31
; 
32'd41231: dataIn1 = 32'd32
; 
32'd41232: dataIn1 = 32'd33
; 
32'd41233: dataIn1 = 32'd34
; 
32'd41234: dataIn1 = 32'd36
; 
32'd41235: dataIn1 = 32'd37
; 
32'd41236: dataIn1 = 32'd38
; 
32'd41237: dataIn1 = 32'd39
; 
32'd41238: dataIn1 = 32'd42
; 
32'd41239: dataIn1 = 32'd44
; 
32'd41240: dataIn1 = 32'd45
; 
32'd41241: dataIn1 = 32'd46
; 
32'd41242: dataIn1 = 32'd47
; 
32'd41243: dataIn1 = 32'd48
; 
32'd41244: dataIn1 = 32'd49
; 
32'd41245: dataIn1 = 32'd50
; 
32'd41246: dataIn1 = 32'd51
; 
32'd41247: dataIn1 = 32'd52
; 
32'd41248: dataIn1 = 32'd53
; 
32'd41249: dataIn1 = 32'd54
; 
32'd41250: dataIn1 = 32'd55
; 
32'd41251: dataIn1 = 32'd56
; 
32'd41252: dataIn1 = 32'd57
; 
32'd41253: dataIn1 = 32'd59
; 
32'd41254: dataIn1 = 32'd60
; 
32'd41255: dataIn1 = 32'd61
; 
32'd41256: dataIn1 = 32'd0
; 
32'd41257: dataIn1 = 32'd1
; 
32'd41258: dataIn1 = 32'd4
; 
32'd41259: dataIn1 = 32'd5
; 
32'd41260: dataIn1 = 32'd6
; 
32'd41261: dataIn1 = 32'd7
; 
32'd41262: dataIn1 = 32'd8
; 
32'd41263: dataIn1 = 32'd9
; 
32'd41264: dataIn1 = 32'd10
; 
32'd41265: dataIn1 = 32'd11
; 
32'd41266: dataIn1 = 32'd12
; 
32'd41267: dataIn1 = 32'd14
; 
32'd41268: dataIn1 = 32'd15
; 
32'd41269: dataIn1 = 32'd16
; 
32'd41270: dataIn1 = 32'd17
; 
32'd41271: dataIn1 = 32'd19
; 
32'd41272: dataIn1 = 32'd20
; 
32'd41273: dataIn1 = 32'd21
; 
32'd41274: dataIn1 = 32'd22
; 
32'd41275: dataIn1 = 32'd23
; 
32'd41276: dataIn1 = 32'd24
; 
32'd41277: dataIn1 = 32'd25
; 
32'd41278: dataIn1 = 32'd26
; 
32'd41279: dataIn1 = 32'd27
; 
32'd41280: dataIn1 = 32'd28
; 
32'd41281: dataIn1 = 32'd29
; 
32'd41282: dataIn1 = 32'd30
; 
32'd41283: dataIn1 = 32'd31
; 
32'd41284: dataIn1 = 32'd32
; 
32'd41285: dataIn1 = 32'd33
; 
32'd41286: dataIn1 = 32'd34
; 
32'd41287: dataIn1 = 32'd35
; 
32'd41288: dataIn1 = 32'd36
; 
32'd41289: dataIn1 = 32'd37
; 
32'd41290: dataIn1 = 32'd38
; 
32'd41291: dataIn1 = 32'd39
; 
32'd41292: dataIn1 = 32'd40
; 
32'd41293: dataIn1 = 32'd42
; 
32'd41294: dataIn1 = 32'd44
; 
32'd41295: dataIn1 = 32'd45
; 
32'd41296: dataIn1 = 32'd47
; 
32'd41297: dataIn1 = 32'd48
; 
32'd41298: dataIn1 = 32'd49
; 
32'd41299: dataIn1 = 32'd50
; 
32'd41300: dataIn1 = 32'd52
; 
32'd41301: dataIn1 = 32'd53
; 
32'd41302: dataIn1 = 32'd54
; 
32'd41303: dataIn1 = 32'd55
; 
32'd41304: dataIn1 = 32'd57
; 
32'd41305: dataIn1 = 32'd58
; 
32'd41306: dataIn1 = 32'd61
; 
32'd41307: dataIn1 = 32'd62
; 
32'd41308: dataIn1 = 32'd63
; 
32'd41309: dataIn1 = 32'd0
; 
32'd41310: dataIn1 = 32'd1
; 
32'd41311: dataIn1 = 32'd2
; 
32'd41312: dataIn1 = 32'd3
; 
32'd41313: dataIn1 = 32'd4
; 
32'd41314: dataIn1 = 32'd5
; 
32'd41315: dataIn1 = 32'd6
; 
32'd41316: dataIn1 = 32'd7
; 
32'd41317: dataIn1 = 32'd8
; 
32'd41318: dataIn1 = 32'd9
; 
32'd41319: dataIn1 = 32'd10
; 
32'd41320: dataIn1 = 32'd11
; 
32'd41321: dataIn1 = 32'd16
; 
32'd41322: dataIn1 = 32'd17
; 
32'd41323: dataIn1 = 32'd18
; 
32'd41324: dataIn1 = 32'd19
; 
32'd41325: dataIn1 = 32'd20
; 
32'd41326: dataIn1 = 32'd21
; 
32'd41327: dataIn1 = 32'd23
; 
32'd41328: dataIn1 = 32'd24
; 
32'd41329: dataIn1 = 32'd25
; 
32'd41330: dataIn1 = 32'd26
; 
32'd41331: dataIn1 = 32'd27
; 
32'd41332: dataIn1 = 32'd29
; 
32'd41333: dataIn1 = 32'd30
; 
32'd41334: dataIn1 = 32'd31
; 
32'd41335: dataIn1 = 32'd32
; 
32'd41336: dataIn1 = 32'd33
; 
32'd41337: dataIn1 = 32'd34
; 
32'd41338: dataIn1 = 32'd35
; 
32'd41339: dataIn1 = 32'd36
; 
32'd41340: dataIn1 = 32'd37
; 
32'd41341: dataIn1 = 32'd38
; 
32'd41342: dataIn1 = 32'd39
; 
32'd41343: dataIn1 = 32'd40
; 
32'd41344: dataIn1 = 32'd42
; 
32'd41345: dataIn1 = 32'd43
; 
32'd41346: dataIn1 = 32'd44
; 
32'd41347: dataIn1 = 32'd45
; 
32'd41348: dataIn1 = 32'd46
; 
32'd41349: dataIn1 = 32'd47
; 
32'd41350: dataIn1 = 32'd48
; 
32'd41351: dataIn1 = 32'd49
; 
32'd41352: dataIn1 = 32'd50
; 
32'd41353: dataIn1 = 32'd51
; 
32'd41354: dataIn1 = 32'd52
; 
32'd41355: dataIn1 = 32'd53
; 
32'd41356: dataIn1 = 32'd54
; 
32'd41357: dataIn1 = 32'd55
; 
32'd41358: dataIn1 = 32'd57
; 
32'd41359: dataIn1 = 32'd58
; 
32'd41360: dataIn1 = 32'd60
; 
32'd41361: dataIn1 = 32'd61
; 
32'd41362: dataIn1 = 32'd62
; 
32'd41363: dataIn1 = 32'd0
; 
32'd41364: dataIn1 = 32'd1
; 
32'd41365: dataIn1 = 32'd2
; 
32'd41366: dataIn1 = 32'd3
; 
32'd41367: dataIn1 = 32'd4
; 
32'd41368: dataIn1 = 32'd5
; 
32'd41369: dataIn1 = 32'd7
; 
32'd41370: dataIn1 = 32'd8
; 
32'd41371: dataIn1 = 32'd9
; 
32'd41372: dataIn1 = 32'd10
; 
32'd41373: dataIn1 = 32'd11
; 
32'd41374: dataIn1 = 32'd12
; 
32'd41375: dataIn1 = 32'd13
; 
32'd41376: dataIn1 = 32'd14
; 
32'd41377: dataIn1 = 32'd15
; 
32'd41378: dataIn1 = 32'd16
; 
32'd41379: dataIn1 = 32'd17
; 
32'd41380: dataIn1 = 32'd18
; 
32'd41381: dataIn1 = 32'd19
; 
32'd41382: dataIn1 = 32'd20
; 
32'd41383: dataIn1 = 32'd21
; 
32'd41384: dataIn1 = 32'd23
; 
32'd41385: dataIn1 = 32'd24
; 
32'd41386: dataIn1 = 32'd25
; 
32'd41387: dataIn1 = 32'd27
; 
32'd41388: dataIn1 = 32'd28
; 
32'd41389: dataIn1 = 32'd30
; 
32'd41390: dataIn1 = 32'd31
; 
32'd41391: dataIn1 = 32'd32
; 
32'd41392: dataIn1 = 32'd33
; 
32'd41393: dataIn1 = 32'd34
; 
32'd41394: dataIn1 = 32'd35
; 
32'd41395: dataIn1 = 32'd36
; 
32'd41396: dataIn1 = 32'd37
; 
32'd41397: dataIn1 = 32'd39
; 
32'd41398: dataIn1 = 32'd40
; 
32'd41399: dataIn1 = 32'd41
; 
32'd41400: dataIn1 = 32'd42
; 
32'd41401: dataIn1 = 32'd43
; 
32'd41402: dataIn1 = 32'd44
; 
32'd41403: dataIn1 = 32'd45
; 
32'd41404: dataIn1 = 32'd47
; 
32'd41405: dataIn1 = 32'd48
; 
32'd41406: dataIn1 = 32'd49
; 
32'd41407: dataIn1 = 32'd51
; 
32'd41408: dataIn1 = 32'd52
; 
32'd41409: dataIn1 = 32'd53
; 
32'd41410: dataIn1 = 32'd54
; 
32'd41411: dataIn1 = 32'd55
; 
32'd41412: dataIn1 = 32'd56
; 
32'd41413: dataIn1 = 32'd57
; 
32'd41414: dataIn1 = 32'd58
; 
32'd41415: dataIn1 = 32'd59
; 
32'd41416: dataIn1 = 32'd60
; 
32'd41417: dataIn1 = 32'd61
; 
32'd41418: dataIn1 = 32'd62
; 
32'd41419: dataIn1 = 32'd63
; 
32'd41420: dataIn1 = 32'd2
; 
32'd41421: dataIn1 = 32'd4
; 
32'd41422: dataIn1 = 32'd5
; 
32'd41423: dataIn1 = 32'd6
; 
32'd41424: dataIn1 = 32'd7
; 
32'd41425: dataIn1 = 32'd9
; 
32'd41426: dataIn1 = 32'd10
; 
32'd41427: dataIn1 = 32'd11
; 
32'd41428: dataIn1 = 32'd12
; 
32'd41429: dataIn1 = 32'd13
; 
32'd41430: dataIn1 = 32'd16
; 
32'd41431: dataIn1 = 32'd17
; 
32'd41432: dataIn1 = 32'd18
; 
32'd41433: dataIn1 = 32'd19
; 
32'd41434: dataIn1 = 32'd20
; 
32'd41435: dataIn1 = 32'd22
; 
32'd41436: dataIn1 = 32'd23
; 
32'd41437: dataIn1 = 32'd24
; 
32'd41438: dataIn1 = 32'd25
; 
32'd41439: dataIn1 = 32'd26
; 
32'd41440: dataIn1 = 32'd27
; 
32'd41441: dataIn1 = 32'd28
; 
32'd41442: dataIn1 = 32'd29
; 
32'd41443: dataIn1 = 32'd30
; 
32'd41444: dataIn1 = 32'd31
; 
32'd41445: dataIn1 = 32'd32
; 
32'd41446: dataIn1 = 32'd33
; 
32'd41447: dataIn1 = 32'd34
; 
32'd41448: dataIn1 = 32'd35
; 
32'd41449: dataIn1 = 32'd36
; 
32'd41450: dataIn1 = 32'd37
; 
32'd41451: dataIn1 = 32'd39
; 
32'd41452: dataIn1 = 32'd40
; 
32'd41453: dataIn1 = 32'd41
; 
32'd41454: dataIn1 = 32'd42
; 
32'd41455: dataIn1 = 32'd43
; 
32'd41456: dataIn1 = 32'd44
; 
32'd41457: dataIn1 = 32'd45
; 
32'd41458: dataIn1 = 32'd46
; 
32'd41459: dataIn1 = 32'd47
; 
32'd41460: dataIn1 = 32'd48
; 
32'd41461: dataIn1 = 32'd49
; 
32'd41462: dataIn1 = 32'd50
; 
32'd41463: dataIn1 = 32'd51
; 
32'd41464: dataIn1 = 32'd52
; 
32'd41465: dataIn1 = 32'd53
; 
32'd41466: dataIn1 = 32'd54
; 
32'd41467: dataIn1 = 32'd55
; 
32'd41468: dataIn1 = 32'd56
; 
32'd41469: dataIn1 = 32'd57
; 
32'd41470: dataIn1 = 32'd58
; 
32'd41471: dataIn1 = 32'd61
; 
32'd41472: dataIn1 = 32'd62
; 
32'd41473: dataIn1 = 32'd63
; 
32'd41474: dataIn1 = 32'd0
; 
32'd41475: dataIn1 = 32'd1
; 
32'd41476: dataIn1 = 32'd2
; 
32'd41477: dataIn1 = 32'd3
; 
32'd41478: dataIn1 = 32'd4
; 
32'd41479: dataIn1 = 32'd5
; 
32'd41480: dataIn1 = 32'd6
; 
32'd41481: dataIn1 = 32'd7
; 
32'd41482: dataIn1 = 32'd9
; 
32'd41483: dataIn1 = 32'd10
; 
32'd41484: dataIn1 = 32'd11
; 
32'd41485: dataIn1 = 32'd12
; 
32'd41486: dataIn1 = 32'd14
; 
32'd41487: dataIn1 = 32'd15
; 
32'd41488: dataIn1 = 32'd16
; 
32'd41489: dataIn1 = 32'd17
; 
32'd41490: dataIn1 = 32'd18
; 
32'd41491: dataIn1 = 32'd20
; 
32'd41492: dataIn1 = 32'd22
; 
32'd41493: dataIn1 = 32'd23
; 
32'd41494: dataIn1 = 32'd24
; 
32'd41495: dataIn1 = 32'd25
; 
32'd41496: dataIn1 = 32'd26
; 
32'd41497: dataIn1 = 32'd27
; 
32'd41498: dataIn1 = 32'd28
; 
32'd41499: dataIn1 = 32'd29
; 
32'd41500: dataIn1 = 32'd30
; 
32'd41501: dataIn1 = 32'd31
; 
32'd41502: dataIn1 = 32'd32
; 
32'd41503: dataIn1 = 32'd33
; 
32'd41504: dataIn1 = 32'd35
; 
32'd41505: dataIn1 = 32'd38
; 
32'd41506: dataIn1 = 32'd39
; 
32'd41507: dataIn1 = 32'd40
; 
32'd41508: dataIn1 = 32'd41
; 
32'd41509: dataIn1 = 32'd43
; 
32'd41510: dataIn1 = 32'd44
; 
32'd41511: dataIn1 = 32'd47
; 
32'd41512: dataIn1 = 32'd49
; 
32'd41513: dataIn1 = 32'd50
; 
32'd41514: dataIn1 = 32'd51
; 
32'd41515: dataIn1 = 32'd53
; 
32'd41516: dataIn1 = 32'd54
; 
32'd41517: dataIn1 = 32'd55
; 
32'd41518: dataIn1 = 32'd56
; 
32'd41519: dataIn1 = 32'd58
; 
32'd41520: dataIn1 = 32'd59
; 
32'd41521: dataIn1 = 32'd60
; 
32'd41522: dataIn1 = 32'd61
; 
32'd41523: dataIn1 = 32'd62
; 
32'd41524: dataIn1 = 32'd63
; 
32'd41525: dataIn1 = 32'd0
; 
32'd41526: dataIn1 = 32'd1
; 
32'd41527: dataIn1 = 32'd3
; 
32'd41528: dataIn1 = 32'd4
; 
32'd41529: dataIn1 = 32'd5
; 
32'd41530: dataIn1 = 32'd7
; 
32'd41531: dataIn1 = 32'd8
; 
32'd41532: dataIn1 = 32'd9
; 
32'd41533: dataIn1 = 32'd10
; 
32'd41534: dataIn1 = 32'd12
; 
32'd41535: dataIn1 = 32'd13
; 
32'd41536: dataIn1 = 32'd14
; 
32'd41537: dataIn1 = 32'd15
; 
32'd41538: dataIn1 = 32'd16
; 
32'd41539: dataIn1 = 32'd17
; 
32'd41540: dataIn1 = 32'd18
; 
32'd41541: dataIn1 = 32'd19
; 
32'd41542: dataIn1 = 32'd20
; 
32'd41543: dataIn1 = 32'd21
; 
32'd41544: dataIn1 = 32'd22
; 
32'd41545: dataIn1 = 32'd23
; 
32'd41546: dataIn1 = 32'd25
; 
32'd41547: dataIn1 = 32'd26
; 
32'd41548: dataIn1 = 32'd27
; 
32'd41549: dataIn1 = 32'd28
; 
32'd41550: dataIn1 = 32'd29
; 
32'd41551: dataIn1 = 32'd30
; 
32'd41552: dataIn1 = 32'd31
; 
32'd41553: dataIn1 = 32'd32
; 
32'd41554: dataIn1 = 32'd33
; 
32'd41555: dataIn1 = 32'd34
; 
32'd41556: dataIn1 = 32'd35
; 
32'd41557: dataIn1 = 32'd37
; 
32'd41558: dataIn1 = 32'd38
; 
32'd41559: dataIn1 = 32'd39
; 
32'd41560: dataIn1 = 32'd40
; 
32'd41561: dataIn1 = 32'd41
; 
32'd41562: dataIn1 = 32'd42
; 
32'd41563: dataIn1 = 32'd43
; 
32'd41564: dataIn1 = 32'd44
; 
32'd41565: dataIn1 = 32'd45
; 
32'd41566: dataIn1 = 32'd46
; 
32'd41567: dataIn1 = 32'd48
; 
32'd41568: dataIn1 = 32'd49
; 
32'd41569: dataIn1 = 32'd51
; 
32'd41570: dataIn1 = 32'd52
; 
32'd41571: dataIn1 = 32'd53
; 
32'd41572: dataIn1 = 32'd55
; 
32'd41573: dataIn1 = 32'd56
; 
32'd41574: dataIn1 = 32'd57
; 
32'd41575: dataIn1 = 32'd58
; 
32'd41576: dataIn1 = 32'd59
; 
32'd41577: dataIn1 = 32'd60
; 
32'd41578: dataIn1 = 32'd61
; 
32'd41579: dataIn1 = 32'd62
; 
32'd41580: dataIn1 = 32'd63
; 
32'd41581: dataIn1 = 32'd0
; 
32'd41582: dataIn1 = 32'd1
; 
32'd41583: dataIn1 = 32'd2
; 
32'd41584: dataIn1 = 32'd3
; 
32'd41585: dataIn1 = 32'd4
; 
32'd41586: dataIn1 = 32'd5
; 
32'd41587: dataIn1 = 32'd6
; 
32'd41588: dataIn1 = 32'd7
; 
32'd41589: dataIn1 = 32'd9
; 
32'd41590: dataIn1 = 32'd10
; 
32'd41591: dataIn1 = 32'd11
; 
32'd41592: dataIn1 = 32'd12
; 
32'd41593: dataIn1 = 32'd13
; 
32'd41594: dataIn1 = 32'd14
; 
32'd41595: dataIn1 = 32'd15
; 
32'd41596: dataIn1 = 32'd16
; 
32'd41597: dataIn1 = 32'd17
; 
32'd41598: dataIn1 = 32'd18
; 
32'd41599: dataIn1 = 32'd19
; 
32'd41600: dataIn1 = 32'd20
; 
32'd41601: dataIn1 = 32'd21
; 
32'd41602: dataIn1 = 32'd22
; 
32'd41603: dataIn1 = 32'd23
; 
32'd41604: dataIn1 = 32'd24
; 
32'd41605: dataIn1 = 32'd25
; 
32'd41606: dataIn1 = 32'd26
; 
32'd41607: dataIn1 = 32'd27
; 
32'd41608: dataIn1 = 32'd28
; 
32'd41609: dataIn1 = 32'd31
; 
32'd41610: dataIn1 = 32'd33
; 
32'd41611: dataIn1 = 32'd34
; 
32'd41612: dataIn1 = 32'd35
; 
32'd41613: dataIn1 = 32'd36
; 
32'd41614: dataIn1 = 32'd37
; 
32'd41615: dataIn1 = 32'd38
; 
32'd41616: dataIn1 = 32'd39
; 
32'd41617: dataIn1 = 32'd40
; 
32'd41618: dataIn1 = 32'd41
; 
32'd41619: dataIn1 = 32'd43
; 
32'd41620: dataIn1 = 32'd44
; 
32'd41621: dataIn1 = 32'd45
; 
32'd41622: dataIn1 = 32'd46
; 
32'd41623: dataIn1 = 32'd47
; 
32'd41624: dataIn1 = 32'd49
; 
32'd41625: dataIn1 = 32'd50
; 
32'd41626: dataIn1 = 32'd51
; 
32'd41627: dataIn1 = 32'd54
; 
32'd41628: dataIn1 = 32'd55
; 
32'd41629: dataIn1 = 32'd56
; 
32'd41630: dataIn1 = 32'd57
; 
32'd41631: dataIn1 = 32'd58
; 
32'd41632: dataIn1 = 32'd59
; 
32'd41633: dataIn1 = 32'd60
; 
32'd41634: dataIn1 = 32'd63
; 
32'd41635: dataIn1 = 32'd0
; 
32'd41636: dataIn1 = 32'd2
; 
32'd41637: dataIn1 = 32'd3
; 
32'd41638: dataIn1 = 32'd4
; 
32'd41639: dataIn1 = 32'd5
; 
32'd41640: dataIn1 = 32'd6
; 
32'd41641: dataIn1 = 32'd7
; 
32'd41642: dataIn1 = 32'd8
; 
32'd41643: dataIn1 = 32'd9
; 
32'd41644: dataIn1 = 32'd10
; 
32'd41645: dataIn1 = 32'd11
; 
32'd41646: dataIn1 = 32'd12
; 
32'd41647: dataIn1 = 32'd13
; 
32'd41648: dataIn1 = 32'd14
; 
32'd41649: dataIn1 = 32'd15
; 
32'd41650: dataIn1 = 32'd16
; 
32'd41651: dataIn1 = 32'd17
; 
32'd41652: dataIn1 = 32'd18
; 
32'd41653: dataIn1 = 32'd19
; 
32'd41654: dataIn1 = 32'd20
; 
32'd41655: dataIn1 = 32'd21
; 
32'd41656: dataIn1 = 32'd22
; 
32'd41657: dataIn1 = 32'd23
; 
32'd41658: dataIn1 = 32'd24
; 
32'd41659: dataIn1 = 32'd25
; 
32'd41660: dataIn1 = 32'd26
; 
32'd41661: dataIn1 = 32'd27
; 
32'd41662: dataIn1 = 32'd28
; 
32'd41663: dataIn1 = 32'd29
; 
32'd41664: dataIn1 = 32'd30
; 
32'd41665: dataIn1 = 32'd31
; 
32'd41666: dataIn1 = 32'd33
; 
32'd41667: dataIn1 = 32'd34
; 
32'd41668: dataIn1 = 32'd35
; 
32'd41669: dataIn1 = 32'd36
; 
32'd41670: dataIn1 = 32'd37
; 
32'd41671: dataIn1 = 32'd38
; 
32'd41672: dataIn1 = 32'd39
; 
32'd41673: dataIn1 = 32'd40
; 
32'd41674: dataIn1 = 32'd41
; 
32'd41675: dataIn1 = 32'd44
; 
32'd41676: dataIn1 = 32'd45
; 
32'd41677: dataIn1 = 32'd46
; 
32'd41678: dataIn1 = 32'd47
; 
32'd41679: dataIn1 = 32'd48
; 
32'd41680: dataIn1 = 32'd49
; 
32'd41681: dataIn1 = 32'd50
; 
32'd41682: dataIn1 = 32'd52
; 
32'd41683: dataIn1 = 32'd53
; 
32'd41684: dataIn1 = 32'd54
; 
32'd41685: dataIn1 = 32'd55
; 
32'd41686: dataIn1 = 32'd56
; 
32'd41687: dataIn1 = 32'd57
; 
32'd41688: dataIn1 = 32'd58
; 
32'd41689: dataIn1 = 32'd59
; 
32'd41690: dataIn1 = 32'd60
; 
32'd41691: dataIn1 = 32'd62
; 
32'd41692: dataIn1 = 32'd63
; 
32'd41693: dataIn1 = 32'd0
; 
32'd41694: dataIn1 = 32'd1
; 
32'd41695: dataIn1 = 32'd2
; 
32'd41696: dataIn1 = 32'd3
; 
32'd41697: dataIn1 = 32'd4
; 
32'd41698: dataIn1 = 32'd5
; 
32'd41699: dataIn1 = 32'd6
; 
32'd41700: dataIn1 = 32'd7
; 
32'd41701: dataIn1 = 32'd8
; 
32'd41702: dataIn1 = 32'd9
; 
32'd41703: dataIn1 = 32'd10
; 
32'd41704: dataIn1 = 32'd11
; 
32'd41705: dataIn1 = 32'd13
; 
32'd41706: dataIn1 = 32'd14
; 
32'd41707: dataIn1 = 32'd15
; 
32'd41708: dataIn1 = 32'd16
; 
32'd41709: dataIn1 = 32'd17
; 
32'd41710: dataIn1 = 32'd18
; 
32'd41711: dataIn1 = 32'd20
; 
32'd41712: dataIn1 = 32'd21
; 
32'd41713: dataIn1 = 32'd22
; 
32'd41714: dataIn1 = 32'd24
; 
32'd41715: dataIn1 = 32'd29
; 
32'd41716: dataIn1 = 32'd30
; 
32'd41717: dataIn1 = 32'd31
; 
32'd41718: dataIn1 = 32'd32
; 
32'd41719: dataIn1 = 32'd33
; 
32'd41720: dataIn1 = 32'd34
; 
32'd41721: dataIn1 = 32'd35
; 
32'd41722: dataIn1 = 32'd36
; 
32'd41723: dataIn1 = 32'd37
; 
32'd41724: dataIn1 = 32'd38
; 
32'd41725: dataIn1 = 32'd39
; 
32'd41726: dataIn1 = 32'd40
; 
32'd41727: dataIn1 = 32'd41
; 
32'd41728: dataIn1 = 32'd43
; 
32'd41729: dataIn1 = 32'd44
; 
32'd41730: dataIn1 = 32'd45
; 
32'd41731: dataIn1 = 32'd46
; 
32'd41732: dataIn1 = 32'd47
; 
32'd41733: dataIn1 = 32'd48
; 
32'd41734: dataIn1 = 32'd49
; 
32'd41735: dataIn1 = 32'd50
; 
32'd41736: dataIn1 = 32'd51
; 
32'd41737: dataIn1 = 32'd52
; 
32'd41738: dataIn1 = 32'd53
; 
32'd41739: dataIn1 = 32'd54
; 
32'd41740: dataIn1 = 32'd55
; 
32'd41741: dataIn1 = 32'd56
; 
32'd41742: dataIn1 = 32'd57
; 
32'd41743: dataIn1 = 32'd59
; 
32'd41744: dataIn1 = 32'd60
; 
32'd41745: dataIn1 = 32'd61
; 
32'd41746: dataIn1 = 32'd63
; 
32'd41747: dataIn1 = 32'd0
; 
32'd41748: dataIn1 = 32'd1
; 
32'd41749: dataIn1 = 32'd2
; 
32'd41750: dataIn1 = 32'd3
; 
32'd41751: dataIn1 = 32'd4
; 
32'd41752: dataIn1 = 32'd5
; 
32'd41753: dataIn1 = 32'd6
; 
32'd41754: dataIn1 = 32'd7
; 
32'd41755: dataIn1 = 32'd8
; 
32'd41756: dataIn1 = 32'd9
; 
32'd41757: dataIn1 = 32'd10
; 
32'd41758: dataIn1 = 32'd11
; 
32'd41759: dataIn1 = 32'd12
; 
32'd41760: dataIn1 = 32'd13
; 
32'd41761: dataIn1 = 32'd14
; 
32'd41762: dataIn1 = 32'd15
; 
32'd41763: dataIn1 = 32'd17
; 
32'd41764: dataIn1 = 32'd18
; 
32'd41765: dataIn1 = 32'd19
; 
32'd41766: dataIn1 = 32'd20
; 
32'd41767: dataIn1 = 32'd21
; 
32'd41768: dataIn1 = 32'd23
; 
32'd41769: dataIn1 = 32'd24
; 
32'd41770: dataIn1 = 32'd25
; 
32'd41771: dataIn1 = 32'd26
; 
32'd41772: dataIn1 = 32'd28
; 
32'd41773: dataIn1 = 32'd29
; 
32'd41774: dataIn1 = 32'd30
; 
32'd41775: dataIn1 = 32'd31
; 
32'd41776: dataIn1 = 32'd32
; 
32'd41777: dataIn1 = 32'd33
; 
32'd41778: dataIn1 = 32'd34
; 
32'd41779: dataIn1 = 32'd35
; 
32'd41780: dataIn1 = 32'd36
; 
32'd41781: dataIn1 = 32'd37
; 
32'd41782: dataIn1 = 32'd38
; 
32'd41783: dataIn1 = 32'd39
; 
32'd41784: dataIn1 = 32'd40
; 
32'd41785: dataIn1 = 32'd41
; 
32'd41786: dataIn1 = 32'd42
; 
32'd41787: dataIn1 = 32'd43
; 
32'd41788: dataIn1 = 32'd44
; 
32'd41789: dataIn1 = 32'd45
; 
32'd41790: dataIn1 = 32'd46
; 
32'd41791: dataIn1 = 32'd47
; 
32'd41792: dataIn1 = 32'd48
; 
32'd41793: dataIn1 = 32'd49
; 
32'd41794: dataIn1 = 32'd50
; 
32'd41795: dataIn1 = 32'd51
; 
32'd41796: dataIn1 = 32'd52
; 
32'd41797: dataIn1 = 32'd53
; 
32'd41798: dataIn1 = 32'd54
; 
32'd41799: dataIn1 = 32'd55
; 
32'd41800: dataIn1 = 32'd56
; 
32'd41801: dataIn1 = 32'd59
; 
32'd41802: dataIn1 = 32'd60
; 
32'd41803: dataIn1 = 32'd61
; 
32'd41804: dataIn1 = 32'd62
; 
32'd41805: dataIn1 = 32'd63
; 
32'd41806: dataIn1 = 32'd0
; 
32'd41807: dataIn1 = 32'd1
; 
32'd41808: dataIn1 = 32'd2
; 
32'd41809: dataIn1 = 32'd3
; 
32'd41810: dataIn1 = 32'd4
; 
32'd41811: dataIn1 = 32'd6
; 
32'd41812: dataIn1 = 32'd7
; 
32'd41813: dataIn1 = 32'd8
; 
32'd41814: dataIn1 = 32'd9
; 
32'd41815: dataIn1 = 32'd11
; 
32'd41816: dataIn1 = 32'd12
; 
32'd41817: dataIn1 = 32'd13
; 
32'd41818: dataIn1 = 32'd15
; 
32'd41819: dataIn1 = 32'd16
; 
32'd41820: dataIn1 = 32'd17
; 
32'd41821: dataIn1 = 32'd18
; 
32'd41822: dataIn1 = 32'd20
; 
32'd41823: dataIn1 = 32'd21
; 
32'd41824: dataIn1 = 32'd22
; 
32'd41825: dataIn1 = 32'd23
; 
32'd41826: dataIn1 = 32'd24
; 
32'd41827: dataIn1 = 32'd25
; 
32'd41828: dataIn1 = 32'd27
; 
32'd41829: dataIn1 = 32'd28
; 
32'd41830: dataIn1 = 32'd29
; 
32'd41831: dataIn1 = 32'd32
; 
32'd41832: dataIn1 = 32'd33
; 
32'd41833: dataIn1 = 32'd34
; 
32'd41834: dataIn1 = 32'd35
; 
32'd41835: dataIn1 = 32'd36
; 
32'd41836: dataIn1 = 32'd37
; 
32'd41837: dataIn1 = 32'd38
; 
32'd41838: dataIn1 = 32'd39
; 
32'd41839: dataIn1 = 32'd40
; 
32'd41840: dataIn1 = 32'd41
; 
32'd41841: dataIn1 = 32'd42
; 
32'd41842: dataIn1 = 32'd43
; 
32'd41843: dataIn1 = 32'd44
; 
32'd41844: dataIn1 = 32'd47
; 
32'd41845: dataIn1 = 32'd48
; 
32'd41846: dataIn1 = 32'd49
; 
32'd41847: dataIn1 = 32'd50
; 
32'd41848: dataIn1 = 32'd51
; 
32'd41849: dataIn1 = 32'd52
; 
32'd41850: dataIn1 = 32'd53
; 
32'd41851: dataIn1 = 32'd54
; 
32'd41852: dataIn1 = 32'd55
; 
32'd41853: dataIn1 = 32'd56
; 
32'd41854: dataIn1 = 32'd57
; 
32'd41855: dataIn1 = 32'd59
; 
32'd41856: dataIn1 = 32'd60
; 
32'd41857: dataIn1 = 32'd61
; 
32'd41858: dataIn1 = 32'd63
; 
32'd41859: dataIn1 = 32'd1
; 
32'd41860: dataIn1 = 32'd2
; 
32'd41861: dataIn1 = 32'd4
; 
32'd41862: dataIn1 = 32'd5
; 
32'd41863: dataIn1 = 32'd6
; 
32'd41864: dataIn1 = 32'd7
; 
32'd41865: dataIn1 = 32'd8
; 
32'd41866: dataIn1 = 32'd9
; 
32'd41867: dataIn1 = 32'd10
; 
32'd41868: dataIn1 = 32'd11
; 
32'd41869: dataIn1 = 32'd12
; 
32'd41870: dataIn1 = 32'd13
; 
32'd41871: dataIn1 = 32'd14
; 
32'd41872: dataIn1 = 32'd15
; 
32'd41873: dataIn1 = 32'd16
; 
32'd41874: dataIn1 = 32'd17
; 
32'd41875: dataIn1 = 32'd18
; 
32'd41876: dataIn1 = 32'd19
; 
32'd41877: dataIn1 = 32'd21
; 
32'd41878: dataIn1 = 32'd22
; 
32'd41879: dataIn1 = 32'd24
; 
32'd41880: dataIn1 = 32'd25
; 
32'd41881: dataIn1 = 32'd26
; 
32'd41882: dataIn1 = 32'd27
; 
32'd41883: dataIn1 = 32'd28
; 
32'd41884: dataIn1 = 32'd29
; 
32'd41885: dataIn1 = 32'd30
; 
32'd41886: dataIn1 = 32'd31
; 
32'd41887: dataIn1 = 32'd32
; 
32'd41888: dataIn1 = 32'd33
; 
32'd41889: dataIn1 = 32'd34
; 
32'd41890: dataIn1 = 32'd35
; 
32'd41891: dataIn1 = 32'd36
; 
32'd41892: dataIn1 = 32'd37
; 
32'd41893: dataIn1 = 32'd38
; 
32'd41894: dataIn1 = 32'd39
; 
32'd41895: dataIn1 = 32'd40
; 
32'd41896: dataIn1 = 32'd41
; 
32'd41897: dataIn1 = 32'd42
; 
32'd41898: dataIn1 = 32'd43
; 
32'd41899: dataIn1 = 32'd44
; 
32'd41900: dataIn1 = 32'd45
; 
32'd41901: dataIn1 = 32'd46
; 
32'd41902: dataIn1 = 32'd47
; 
32'd41903: dataIn1 = 32'd49
; 
32'd41904: dataIn1 = 32'd50
; 
32'd41905: dataIn1 = 32'd52
; 
32'd41906: dataIn1 = 32'd53
; 
32'd41907: dataIn1 = 32'd54
; 
32'd41908: dataIn1 = 32'd55
; 
32'd41909: dataIn1 = 32'd56
; 
32'd41910: dataIn1 = 32'd57
; 
32'd41911: dataIn1 = 32'd59
; 
32'd41912: dataIn1 = 32'd61
; 
32'd41913: dataIn1 = 32'd62
; 
32'd41914: dataIn1 = 32'd1
; 
32'd41915: dataIn1 = 32'd2
; 
32'd41916: dataIn1 = 32'd6
; 
32'd41917: dataIn1 = 32'd7
; 
32'd41918: dataIn1 = 32'd8
; 
32'd41919: dataIn1 = 32'd9
; 
32'd41920: dataIn1 = 32'd10
; 
32'd41921: dataIn1 = 32'd11
; 
32'd41922: dataIn1 = 32'd12
; 
32'd41923: dataIn1 = 32'd15
; 
32'd41924: dataIn1 = 32'd16
; 
32'd41925: dataIn1 = 32'd17
; 
32'd41926: dataIn1 = 32'd18
; 
32'd41927: dataIn1 = 32'd19
; 
32'd41928: dataIn1 = 32'd20
; 
32'd41929: dataIn1 = 32'd21
; 
32'd41930: dataIn1 = 32'd23
; 
32'd41931: dataIn1 = 32'd24
; 
32'd41932: dataIn1 = 32'd25
; 
32'd41933: dataIn1 = 32'd26
; 
32'd41934: dataIn1 = 32'd27
; 
32'd41935: dataIn1 = 32'd30
; 
32'd41936: dataIn1 = 32'd31
; 
32'd41937: dataIn1 = 32'd32
; 
32'd41938: dataIn1 = 32'd33
; 
32'd41939: dataIn1 = 32'd34
; 
32'd41940: dataIn1 = 32'd35
; 
32'd41941: dataIn1 = 32'd36
; 
32'd41942: dataIn1 = 32'd38
; 
32'd41943: dataIn1 = 32'd40
; 
32'd41944: dataIn1 = 32'd41
; 
32'd41945: dataIn1 = 32'd42
; 
32'd41946: dataIn1 = 32'd45
; 
32'd41947: dataIn1 = 32'd46
; 
32'd41948: dataIn1 = 32'd47
; 
32'd41949: dataIn1 = 32'd48
; 
32'd41950: dataIn1 = 32'd49
; 
32'd41951: dataIn1 = 32'd51
; 
32'd41952: dataIn1 = 32'd53
; 
32'd41953: dataIn1 = 32'd54
; 
32'd41954: dataIn1 = 32'd55
; 
32'd41955: dataIn1 = 32'd56
; 
32'd41956: dataIn1 = 32'd57
; 
32'd41957: dataIn1 = 32'd58
; 
32'd41958: dataIn1 = 32'd59
; 
32'd41959: dataIn1 = 32'd60
; 
32'd41960: dataIn1 = 32'd61
; 
32'd41961: dataIn1 = 32'd62
; 
32'd41962: dataIn1 = 32'd63
; 
32'd41963: dataIn1 = 32'd0
; 
32'd41964: dataIn1 = 32'd1
; 
32'd41965: dataIn1 = 32'd2
; 
32'd41966: dataIn1 = 32'd3
; 
32'd41967: dataIn1 = 32'd4
; 
32'd41968: dataIn1 = 32'd5
; 
32'd41969: dataIn1 = 32'd6
; 
32'd41970: dataIn1 = 32'd8
; 
32'd41971: dataIn1 = 32'd9
; 
32'd41972: dataIn1 = 32'd10
; 
32'd41973: dataIn1 = 32'd11
; 
32'd41974: dataIn1 = 32'd12
; 
32'd41975: dataIn1 = 32'd13
; 
32'd41976: dataIn1 = 32'd14
; 
32'd41977: dataIn1 = 32'd15
; 
32'd41978: dataIn1 = 32'd17
; 
32'd41979: dataIn1 = 32'd19
; 
32'd41980: dataIn1 = 32'd20
; 
32'd41981: dataIn1 = 32'd21
; 
32'd41982: dataIn1 = 32'd22
; 
32'd41983: dataIn1 = 32'd23
; 
32'd41984: dataIn1 = 32'd24
; 
32'd41985: dataIn1 = 32'd25
; 
32'd41986: dataIn1 = 32'd26
; 
32'd41987: dataIn1 = 32'd27
; 
32'd41988: dataIn1 = 32'd29
; 
32'd41989: dataIn1 = 32'd30
; 
32'd41990: dataIn1 = 32'd31
; 
32'd41991: dataIn1 = 32'd33
; 
32'd41992: dataIn1 = 32'd34
; 
32'd41993: dataIn1 = 32'd35
; 
32'd41994: dataIn1 = 32'd37
; 
32'd41995: dataIn1 = 32'd38
; 
32'd41996: dataIn1 = 32'd39
; 
32'd41997: dataIn1 = 32'd40
; 
32'd41998: dataIn1 = 32'd41
; 
32'd41999: dataIn1 = 32'd42
; 
32'd42000: dataIn1 = 32'd43
; 
32'd42001: dataIn1 = 32'd44
; 
32'd42002: dataIn1 = 32'd45
; 
32'd42003: dataIn1 = 32'd47
; 
32'd42004: dataIn1 = 32'd48
; 
32'd42005: dataIn1 = 32'd50
; 
32'd42006: dataIn1 = 32'd52
; 
32'd42007: dataIn1 = 32'd53
; 
32'd42008: dataIn1 = 32'd54
; 
32'd42009: dataIn1 = 32'd55
; 
32'd42010: dataIn1 = 32'd56
; 
32'd42011: dataIn1 = 32'd57
; 
32'd42012: dataIn1 = 32'd58
; 
32'd42013: dataIn1 = 32'd59
; 
32'd42014: dataIn1 = 32'd60
; 
32'd42015: dataIn1 = 32'd61
; 
32'd42016: dataIn1 = 32'd62
; 
32'd42017: dataIn1 = 32'd63
; 
32'd42018: dataIn1 = 32'd0
; 
32'd42019: dataIn1 = 32'd1
; 
32'd42020: dataIn1 = 32'd2
; 
32'd42021: dataIn1 = 32'd3
; 
32'd42022: dataIn1 = 32'd4
; 
32'd42023: dataIn1 = 32'd5
; 
32'd42024: dataIn1 = 32'd6
; 
32'd42025: dataIn1 = 32'd7
; 
32'd42026: dataIn1 = 32'd8
; 
32'd42027: dataIn1 = 32'd10
; 
32'd42028: dataIn1 = 32'd11
; 
32'd42029: dataIn1 = 32'd12
; 
32'd42030: dataIn1 = 32'd13
; 
32'd42031: dataIn1 = 32'd14
; 
32'd42032: dataIn1 = 32'd15
; 
32'd42033: dataIn1 = 32'd16
; 
32'd42034: dataIn1 = 32'd17
; 
32'd42035: dataIn1 = 32'd18
; 
32'd42036: dataIn1 = 32'd19
; 
32'd42037: dataIn1 = 32'd20
; 
32'd42038: dataIn1 = 32'd22
; 
32'd42039: dataIn1 = 32'd23
; 
32'd42040: dataIn1 = 32'd24
; 
32'd42041: dataIn1 = 32'd25
; 
32'd42042: dataIn1 = 32'd28
; 
32'd42043: dataIn1 = 32'd30
; 
32'd42044: dataIn1 = 32'd31
; 
32'd42045: dataIn1 = 32'd32
; 
32'd42046: dataIn1 = 32'd33
; 
32'd42047: dataIn1 = 32'd34
; 
32'd42048: dataIn1 = 32'd35
; 
32'd42049: dataIn1 = 32'd36
; 
32'd42050: dataIn1 = 32'd37
; 
32'd42051: dataIn1 = 32'd41
; 
32'd42052: dataIn1 = 32'd42
; 
32'd42053: dataIn1 = 32'd43
; 
32'd42054: dataIn1 = 32'd44
; 
32'd42055: dataIn1 = 32'd48
; 
32'd42056: dataIn1 = 32'd49
; 
32'd42057: dataIn1 = 32'd50
; 
32'd42058: dataIn1 = 32'd52
; 
32'd42059: dataIn1 = 32'd53
; 
32'd42060: dataIn1 = 32'd54
; 
32'd42061: dataIn1 = 32'd56
; 
32'd42062: dataIn1 = 32'd57
; 
32'd42063: dataIn1 = 32'd58
; 
32'd42064: dataIn1 = 32'd59
; 
32'd42065: dataIn1 = 32'd60
; 
32'd42066: dataIn1 = 32'd62
; 
32'd42067: dataIn1 = 32'd63
; 
32'd42068: dataIn1 = 32'd0
; 
32'd42069: dataIn1 = 32'd1
; 
32'd42070: dataIn1 = 32'd2
; 
32'd42071: dataIn1 = 32'd3
; 
32'd42072: dataIn1 = 32'd4
; 
32'd42073: dataIn1 = 32'd6
; 
32'd42074: dataIn1 = 32'd8
; 
32'd42075: dataIn1 = 32'd9
; 
32'd42076: dataIn1 = 32'd10
; 
32'd42077: dataIn1 = 32'd11
; 
32'd42078: dataIn1 = 32'd12
; 
32'd42079: dataIn1 = 32'd13
; 
32'd42080: dataIn1 = 32'd14
; 
32'd42081: dataIn1 = 32'd15
; 
32'd42082: dataIn1 = 32'd18
; 
32'd42083: dataIn1 = 32'd19
; 
32'd42084: dataIn1 = 32'd20
; 
32'd42085: dataIn1 = 32'd21
; 
32'd42086: dataIn1 = 32'd22
; 
32'd42087: dataIn1 = 32'd23
; 
32'd42088: dataIn1 = 32'd24
; 
32'd42089: dataIn1 = 32'd25
; 
32'd42090: dataIn1 = 32'd26
; 
32'd42091: dataIn1 = 32'd28
; 
32'd42092: dataIn1 = 32'd29
; 
32'd42093: dataIn1 = 32'd30
; 
32'd42094: dataIn1 = 32'd32
; 
32'd42095: dataIn1 = 32'd33
; 
32'd42096: dataIn1 = 32'd34
; 
32'd42097: dataIn1 = 32'd35
; 
32'd42098: dataIn1 = 32'd36
; 
32'd42099: dataIn1 = 32'd37
; 
32'd42100: dataIn1 = 32'd38
; 
32'd42101: dataIn1 = 32'd39
; 
32'd42102: dataIn1 = 32'd40
; 
32'd42103: dataIn1 = 32'd41
; 
32'd42104: dataIn1 = 32'd42
; 
32'd42105: dataIn1 = 32'd43
; 
32'd42106: dataIn1 = 32'd44
; 
32'd42107: dataIn1 = 32'd45
; 
32'd42108: dataIn1 = 32'd47
; 
32'd42109: dataIn1 = 32'd48
; 
32'd42110: dataIn1 = 32'd49
; 
32'd42111: dataIn1 = 32'd50
; 
32'd42112: dataIn1 = 32'd51
; 
32'd42113: dataIn1 = 32'd52
; 
32'd42114: dataIn1 = 32'd53
; 
32'd42115: dataIn1 = 32'd54
; 
32'd42116: dataIn1 = 32'd57
; 
32'd42117: dataIn1 = 32'd58
; 
32'd42118: dataIn1 = 32'd59
; 
32'd42119: dataIn1 = 32'd60
; 
32'd42120: dataIn1 = 32'd61
; 
32'd42121: dataIn1 = 32'd62
; 
32'd42122: dataIn1 = 32'd63
; 
32'd42123: dataIn1 = 32'd0
; 
32'd42124: dataIn1 = 32'd1
; 
32'd42125: dataIn1 = 32'd2
; 
32'd42126: dataIn1 = 32'd3
; 
32'd42127: dataIn1 = 32'd4
; 
32'd42128: dataIn1 = 32'd5
; 
32'd42129: dataIn1 = 32'd6
; 
32'd42130: dataIn1 = 32'd7
; 
32'd42131: dataIn1 = 32'd8
; 
32'd42132: dataIn1 = 32'd9
; 
32'd42133: dataIn1 = 32'd10
; 
32'd42134: dataIn1 = 32'd11
; 
32'd42135: dataIn1 = 32'd13
; 
32'd42136: dataIn1 = 32'd15
; 
32'd42137: dataIn1 = 32'd17
; 
32'd42138: dataIn1 = 32'd18
; 
32'd42139: dataIn1 = 32'd20
; 
32'd42140: dataIn1 = 32'd21
; 
32'd42141: dataIn1 = 32'd22
; 
32'd42142: dataIn1 = 32'd23
; 
32'd42143: dataIn1 = 32'd24
; 
32'd42144: dataIn1 = 32'd25
; 
32'd42145: dataIn1 = 32'd26
; 
32'd42146: dataIn1 = 32'd27
; 
32'd42147: dataIn1 = 32'd29
; 
32'd42148: dataIn1 = 32'd30
; 
32'd42149: dataIn1 = 32'd31
; 
32'd42150: dataIn1 = 32'd32
; 
32'd42151: dataIn1 = 32'd33
; 
32'd42152: dataIn1 = 32'd34
; 
32'd42153: dataIn1 = 32'd35
; 
32'd42154: dataIn1 = 32'd36
; 
32'd42155: dataIn1 = 32'd38
; 
32'd42156: dataIn1 = 32'd39
; 
32'd42157: dataIn1 = 32'd40
; 
32'd42158: dataIn1 = 32'd42
; 
32'd42159: dataIn1 = 32'd43
; 
32'd42160: dataIn1 = 32'd44
; 
32'd42161: dataIn1 = 32'd45
; 
32'd42162: dataIn1 = 32'd46
; 
32'd42163: dataIn1 = 32'd47
; 
32'd42164: dataIn1 = 32'd48
; 
32'd42165: dataIn1 = 32'd49
; 
32'd42166: dataIn1 = 32'd50
; 
32'd42167: dataIn1 = 32'd52
; 
32'd42168: dataIn1 = 32'd53
; 
32'd42169: dataIn1 = 32'd54
; 
32'd42170: dataIn1 = 32'd55
; 
32'd42171: dataIn1 = 32'd56
; 
32'd42172: dataIn1 = 32'd57
; 
32'd42173: dataIn1 = 32'd58
; 
32'd42174: dataIn1 = 32'd59
; 
32'd42175: dataIn1 = 32'd60
; 
32'd42176: dataIn1 = 32'd61
; 
32'd42177: dataIn1 = 32'd62
; 
32'd42178: dataIn1 = 32'd63
; 
32'd42179: dataIn1 = 32'd0
; 
32'd42180: dataIn1 = 32'd1
; 
32'd42181: dataIn1 = 32'd2
; 
32'd42182: dataIn1 = 32'd3
; 
32'd42183: dataIn1 = 32'd4
; 
32'd42184: dataIn1 = 32'd5
; 
32'd42185: dataIn1 = 32'd6
; 
32'd42186: dataIn1 = 32'd7
; 
32'd42187: dataIn1 = 32'd8
; 
32'd42188: dataIn1 = 32'd9
; 
32'd42189: dataIn1 = 32'd10
; 
32'd42190: dataIn1 = 32'd12
; 
32'd42191: dataIn1 = 32'd13
; 
32'd42192: dataIn1 = 32'd14
; 
32'd42193: dataIn1 = 32'd15
; 
32'd42194: dataIn1 = 32'd16
; 
32'd42195: dataIn1 = 32'd17
; 
32'd42196: dataIn1 = 32'd18
; 
32'd42197: dataIn1 = 32'd19
; 
32'd42198: dataIn1 = 32'd20
; 
32'd42199: dataIn1 = 32'd21
; 
32'd42200: dataIn1 = 32'd22
; 
32'd42201: dataIn1 = 32'd23
; 
32'd42202: dataIn1 = 32'd24
; 
32'd42203: dataIn1 = 32'd25
; 
32'd42204: dataIn1 = 32'd26
; 
32'd42205: dataIn1 = 32'd27
; 
32'd42206: dataIn1 = 32'd29
; 
32'd42207: dataIn1 = 32'd30
; 
32'd42208: dataIn1 = 32'd31
; 
32'd42209: dataIn1 = 32'd33
; 
32'd42210: dataIn1 = 32'd34
; 
32'd42211: dataIn1 = 32'd35
; 
32'd42212: dataIn1 = 32'd36
; 
32'd42213: dataIn1 = 32'd37
; 
32'd42214: dataIn1 = 32'd38
; 
32'd42215: dataIn1 = 32'd39
; 
32'd42216: dataIn1 = 32'd40
; 
32'd42217: dataIn1 = 32'd41
; 
32'd42218: dataIn1 = 32'd42
; 
32'd42219: dataIn1 = 32'd43
; 
32'd42220: dataIn1 = 32'd44
; 
32'd42221: dataIn1 = 32'd45
; 
32'd42222: dataIn1 = 32'd46
; 
32'd42223: dataIn1 = 32'd47
; 
32'd42224: dataIn1 = 32'd50
; 
32'd42225: dataIn1 = 32'd51
; 
32'd42226: dataIn1 = 32'd52
; 
32'd42227: dataIn1 = 32'd53
; 
32'd42228: dataIn1 = 32'd54
; 
32'd42229: dataIn1 = 32'd55
; 
32'd42230: dataIn1 = 32'd56
; 
32'd42231: dataIn1 = 32'd57
; 
32'd42232: dataIn1 = 32'd58
; 
32'd42233: dataIn1 = 32'd59
; 
32'd42234: dataIn1 = 32'd61
; 
32'd42235: dataIn1 = 32'd62
; 
32'd42236: dataIn1 = 32'd63
; 
32'd42237: dataIn1 = 32'd0
; 
32'd42238: dataIn1 = 32'd1
; 
32'd42239: dataIn1 = 32'd3
; 
32'd42240: dataIn1 = 32'd5
; 
32'd42241: dataIn1 = 32'd6
; 
32'd42242: dataIn1 = 32'd8
; 
32'd42243: dataIn1 = 32'd9
; 
32'd42244: dataIn1 = 32'd10
; 
32'd42245: dataIn1 = 32'd11
; 
32'd42246: dataIn1 = 32'd12
; 
32'd42247: dataIn1 = 32'd13
; 
32'd42248: dataIn1 = 32'd14
; 
32'd42249: dataIn1 = 32'd15
; 
32'd42250: dataIn1 = 32'd16
; 
32'd42251: dataIn1 = 32'd17
; 
32'd42252: dataIn1 = 32'd18
; 
32'd42253: dataIn1 = 32'd19
; 
32'd42254: dataIn1 = 32'd20
; 
32'd42255: dataIn1 = 32'd21
; 
32'd42256: dataIn1 = 32'd23
; 
32'd42257: dataIn1 = 32'd24
; 
32'd42258: dataIn1 = 32'd25
; 
32'd42259: dataIn1 = 32'd26
; 
32'd42260: dataIn1 = 32'd27
; 
32'd42261: dataIn1 = 32'd29
; 
32'd42262: dataIn1 = 32'd30
; 
32'd42263: dataIn1 = 32'd31
; 
32'd42264: dataIn1 = 32'd32
; 
32'd42265: dataIn1 = 32'd33
; 
32'd42266: dataIn1 = 32'd34
; 
32'd42267: dataIn1 = 32'd35
; 
32'd42268: dataIn1 = 32'd36
; 
32'd42269: dataIn1 = 32'd37
; 
32'd42270: dataIn1 = 32'd38
; 
32'd42271: dataIn1 = 32'd39
; 
32'd42272: dataIn1 = 32'd41
; 
32'd42273: dataIn1 = 32'd42
; 
32'd42274: dataIn1 = 32'd44
; 
32'd42275: dataIn1 = 32'd45
; 
32'd42276: dataIn1 = 32'd47
; 
32'd42277: dataIn1 = 32'd48
; 
32'd42278: dataIn1 = 32'd49
; 
32'd42279: dataIn1 = 32'd50
; 
32'd42280: dataIn1 = 32'd51
; 
32'd42281: dataIn1 = 32'd52
; 
32'd42282: dataIn1 = 32'd53
; 
32'd42283: dataIn1 = 32'd54
; 
32'd42284: dataIn1 = 32'd55
; 
32'd42285: dataIn1 = 32'd56
; 
32'd42286: dataIn1 = 32'd57
; 
32'd42287: dataIn1 = 32'd58
; 
32'd42288: dataIn1 = 32'd59
; 
32'd42289: dataIn1 = 32'd61
; 
32'd42290: dataIn1 = 32'd62
; 
32'd42291: dataIn1 = 32'd63
; 
32'd42292: dataIn1 = 32'd0
; 
32'd42293: dataIn1 = 32'd1
; 
32'd42294: dataIn1 = 32'd2
; 
32'd42295: dataIn1 = 32'd3
; 
32'd42296: dataIn1 = 32'd4
; 
32'd42297: dataIn1 = 32'd5
; 
32'd42298: dataIn1 = 32'd6
; 
32'd42299: dataIn1 = 32'd8
; 
32'd42300: dataIn1 = 32'd9
; 
32'd42301: dataIn1 = 32'd10
; 
32'd42302: dataIn1 = 32'd11
; 
32'd42303: dataIn1 = 32'd13
; 
32'd42304: dataIn1 = 32'd14
; 
32'd42305: dataIn1 = 32'd15
; 
32'd42306: dataIn1 = 32'd16
; 
32'd42307: dataIn1 = 32'd18
; 
32'd42308: dataIn1 = 32'd19
; 
32'd42309: dataIn1 = 32'd20
; 
32'd42310: dataIn1 = 32'd21
; 
32'd42311: dataIn1 = 32'd22
; 
32'd42312: dataIn1 = 32'd23
; 
32'd42313: dataIn1 = 32'd24
; 
32'd42314: dataIn1 = 32'd25
; 
32'd42315: dataIn1 = 32'd26
; 
32'd42316: dataIn1 = 32'd28
; 
32'd42317: dataIn1 = 32'd29
; 
32'd42318: dataIn1 = 32'd31
; 
32'd42319: dataIn1 = 32'd32
; 
32'd42320: dataIn1 = 32'd33
; 
32'd42321: dataIn1 = 32'd35
; 
32'd42322: dataIn1 = 32'd36
; 
32'd42323: dataIn1 = 32'd37
; 
32'd42324: dataIn1 = 32'd38
; 
32'd42325: dataIn1 = 32'd39
; 
32'd42326: dataIn1 = 32'd40
; 
32'd42327: dataIn1 = 32'd42
; 
32'd42328: dataIn1 = 32'd43
; 
32'd42329: dataIn1 = 32'd44
; 
32'd42330: dataIn1 = 32'd45
; 
32'd42331: dataIn1 = 32'd46
; 
32'd42332: dataIn1 = 32'd47
; 
32'd42333: dataIn1 = 32'd48
; 
32'd42334: dataIn1 = 32'd49
; 
32'd42335: dataIn1 = 32'd51
; 
32'd42336: dataIn1 = 32'd53
; 
32'd42337: dataIn1 = 32'd54
; 
32'd42338: dataIn1 = 32'd57
; 
32'd42339: dataIn1 = 32'd59
; 
32'd42340: dataIn1 = 32'd60
; 
32'd42341: dataIn1 = 32'd0
; 
32'd42342: dataIn1 = 32'd1
; 
32'd42343: dataIn1 = 32'd2
; 
32'd42344: dataIn1 = 32'd4
; 
32'd42345: dataIn1 = 32'd5
; 
32'd42346: dataIn1 = 32'd6
; 
32'd42347: dataIn1 = 32'd7
; 
32'd42348: dataIn1 = 32'd9
; 
32'd42349: dataIn1 = 32'd11
; 
32'd42350: dataIn1 = 32'd12
; 
32'd42351: dataIn1 = 32'd13
; 
32'd42352: dataIn1 = 32'd14
; 
32'd42353: dataIn1 = 32'd15
; 
32'd42354: dataIn1 = 32'd16
; 
32'd42355: dataIn1 = 32'd18
; 
32'd42356: dataIn1 = 32'd19
; 
32'd42357: dataIn1 = 32'd20
; 
32'd42358: dataIn1 = 32'd21
; 
32'd42359: dataIn1 = 32'd22
; 
32'd42360: dataIn1 = 32'd23
; 
32'd42361: dataIn1 = 32'd24
; 
32'd42362: dataIn1 = 32'd25
; 
32'd42363: dataIn1 = 32'd26
; 
32'd42364: dataIn1 = 32'd27
; 
32'd42365: dataIn1 = 32'd28
; 
32'd42366: dataIn1 = 32'd29
; 
32'd42367: dataIn1 = 32'd30
; 
32'd42368: dataIn1 = 32'd31
; 
32'd42369: dataIn1 = 32'd32
; 
32'd42370: dataIn1 = 32'd33
; 
32'd42371: dataIn1 = 32'd34
; 
32'd42372: dataIn1 = 32'd35
; 
32'd42373: dataIn1 = 32'd36
; 
32'd42374: dataIn1 = 32'd38
; 
32'd42375: dataIn1 = 32'd39
; 
32'd42376: dataIn1 = 32'd40
; 
32'd42377: dataIn1 = 32'd41
; 
32'd42378: dataIn1 = 32'd42
; 
32'd42379: dataIn1 = 32'd43
; 
32'd42380: dataIn1 = 32'd44
; 
32'd42381: dataIn1 = 32'd45
; 
32'd42382: dataIn1 = 32'd46
; 
32'd42383: dataIn1 = 32'd47
; 
32'd42384: dataIn1 = 32'd48
; 
32'd42385: dataIn1 = 32'd49
; 
32'd42386: dataIn1 = 32'd50
; 
32'd42387: dataIn1 = 32'd51
; 
32'd42388: dataIn1 = 32'd52
; 
32'd42389: dataIn1 = 32'd53
; 
32'd42390: dataIn1 = 32'd54
; 
32'd42391: dataIn1 = 32'd55
; 
32'd42392: dataIn1 = 32'd57
; 
32'd42393: dataIn1 = 32'd58
; 
32'd42394: dataIn1 = 32'd59
; 
32'd42395: dataIn1 = 32'd60
; 
32'd42396: dataIn1 = 32'd61
; 
32'd42397: dataIn1 = 32'd63
; 
32'd42398: dataIn1 = 32'd0
; 
32'd42399: dataIn1 = 32'd1
; 
32'd42400: dataIn1 = 32'd2
; 
32'd42401: dataIn1 = 32'd4
; 
32'd42402: dataIn1 = 32'd5
; 
32'd42403: dataIn1 = 32'd6
; 
32'd42404: dataIn1 = 32'd7
; 
32'd42405: dataIn1 = 32'd8
; 
32'd42406: dataIn1 = 32'd10
; 
32'd42407: dataIn1 = 32'd11
; 
32'd42408: dataIn1 = 32'd12
; 
32'd42409: dataIn1 = 32'd14
; 
32'd42410: dataIn1 = 32'd15
; 
32'd42411: dataIn1 = 32'd16
; 
32'd42412: dataIn1 = 32'd17
; 
32'd42413: dataIn1 = 32'd18
; 
32'd42414: dataIn1 = 32'd19
; 
32'd42415: dataIn1 = 32'd20
; 
32'd42416: dataIn1 = 32'd21
; 
32'd42417: dataIn1 = 32'd23
; 
32'd42418: dataIn1 = 32'd24
; 
32'd42419: dataIn1 = 32'd25
; 
32'd42420: dataIn1 = 32'd26
; 
32'd42421: dataIn1 = 32'd27
; 
32'd42422: dataIn1 = 32'd28
; 
32'd42423: dataIn1 = 32'd29
; 
32'd42424: dataIn1 = 32'd30
; 
32'd42425: dataIn1 = 32'd32
; 
32'd42426: dataIn1 = 32'd33
; 
32'd42427: dataIn1 = 32'd34
; 
32'd42428: dataIn1 = 32'd35
; 
32'd42429: dataIn1 = 32'd37
; 
32'd42430: dataIn1 = 32'd38
; 
32'd42431: dataIn1 = 32'd39
; 
32'd42432: dataIn1 = 32'd40
; 
32'd42433: dataIn1 = 32'd41
; 
32'd42434: dataIn1 = 32'd42
; 
32'd42435: dataIn1 = 32'd43
; 
32'd42436: dataIn1 = 32'd44
; 
32'd42437: dataIn1 = 32'd45
; 
32'd42438: dataIn1 = 32'd46
; 
32'd42439: dataIn1 = 32'd47
; 
32'd42440: dataIn1 = 32'd48
; 
32'd42441: dataIn1 = 32'd49
; 
32'd42442: dataIn1 = 32'd50
; 
32'd42443: dataIn1 = 32'd51
; 
32'd42444: dataIn1 = 32'd52
; 
32'd42445: dataIn1 = 32'd53
; 
32'd42446: dataIn1 = 32'd54
; 
32'd42447: dataIn1 = 32'd55
; 
32'd42448: dataIn1 = 32'd56
; 
32'd42449: dataIn1 = 32'd58
; 
32'd42450: dataIn1 = 32'd59
; 
32'd42451: dataIn1 = 32'd60
; 
32'd42452: dataIn1 = 32'd61
; 
32'd42453: dataIn1 = 32'd62
; 
32'd42454: dataIn1 = 32'd63
; 
32'd42455: dataIn1 = 32'd0
; 
32'd42456: dataIn1 = 32'd1
; 
32'd42457: dataIn1 = 32'd2
; 
32'd42458: dataIn1 = 32'd3
; 
32'd42459: dataIn1 = 32'd4
; 
32'd42460: dataIn1 = 32'd5
; 
32'd42461: dataIn1 = 32'd6
; 
32'd42462: dataIn1 = 32'd8
; 
32'd42463: dataIn1 = 32'd9
; 
32'd42464: dataIn1 = 32'd11
; 
32'd42465: dataIn1 = 32'd12
; 
32'd42466: dataIn1 = 32'd13
; 
32'd42467: dataIn1 = 32'd14
; 
32'd42468: dataIn1 = 32'd15
; 
32'd42469: dataIn1 = 32'd16
; 
32'd42470: dataIn1 = 32'd17
; 
32'd42471: dataIn1 = 32'd18
; 
32'd42472: dataIn1 = 32'd19
; 
32'd42473: dataIn1 = 32'd20
; 
32'd42474: dataIn1 = 32'd21
; 
32'd42475: dataIn1 = 32'd22
; 
32'd42476: dataIn1 = 32'd23
; 
32'd42477: dataIn1 = 32'd24
; 
32'd42478: dataIn1 = 32'd25
; 
32'd42479: dataIn1 = 32'd26
; 
32'd42480: dataIn1 = 32'd27
; 
32'd42481: dataIn1 = 32'd28
; 
32'd42482: dataIn1 = 32'd29
; 
32'd42483: dataIn1 = 32'd30
; 
32'd42484: dataIn1 = 32'd31
; 
32'd42485: dataIn1 = 32'd32
; 
32'd42486: dataIn1 = 32'd33
; 
32'd42487: dataIn1 = 32'd34
; 
32'd42488: dataIn1 = 32'd35
; 
32'd42489: dataIn1 = 32'd36
; 
32'd42490: dataIn1 = 32'd37
; 
32'd42491: dataIn1 = 32'd38
; 
32'd42492: dataIn1 = 32'd39
; 
32'd42493: dataIn1 = 32'd40
; 
32'd42494: dataIn1 = 32'd42
; 
32'd42495: dataIn1 = 32'd43
; 
32'd42496: dataIn1 = 32'd44
; 
32'd42497: dataIn1 = 32'd45
; 
32'd42498: dataIn1 = 32'd46
; 
32'd42499: dataIn1 = 32'd47
; 
32'd42500: dataIn1 = 32'd48
; 
32'd42501: dataIn1 = 32'd49
; 
32'd42502: dataIn1 = 32'd51
; 
32'd42503: dataIn1 = 32'd52
; 
32'd42504: dataIn1 = 32'd53
; 
32'd42505: dataIn1 = 32'd54
; 
32'd42506: dataIn1 = 32'd55
; 
32'd42507: dataIn1 = 32'd56
; 
32'd42508: dataIn1 = 32'd57
; 
32'd42509: dataIn1 = 32'd58
; 
32'd42510: dataIn1 = 32'd59
; 
32'd42511: dataIn1 = 32'd60
; 
32'd42512: dataIn1 = 32'd61
; 
32'd42513: dataIn1 = 32'd62
; 
32'd42514: dataIn1 = 32'd63
; 
32'd42515: dataIn1 = 32'd0
; 
32'd42516: dataIn1 = 32'd1
; 
32'd42517: dataIn1 = 32'd2
; 
32'd42518: dataIn1 = 32'd3
; 
32'd42519: dataIn1 = 32'd4
; 
32'd42520: dataIn1 = 32'd5
; 
32'd42521: dataIn1 = 32'd6
; 
32'd42522: dataIn1 = 32'd7
; 
32'd42523: dataIn1 = 32'd8
; 
32'd42524: dataIn1 = 32'd9
; 
32'd42525: dataIn1 = 32'd10
; 
32'd42526: dataIn1 = 32'd11
; 
32'd42527: dataIn1 = 32'd12
; 
32'd42528: dataIn1 = 32'd13
; 
32'd42529: dataIn1 = 32'd14
; 
32'd42530: dataIn1 = 32'd15
; 
32'd42531: dataIn1 = 32'd16
; 
32'd42532: dataIn1 = 32'd18
; 
32'd42533: dataIn1 = 32'd19
; 
32'd42534: dataIn1 = 32'd21
; 
32'd42535: dataIn1 = 32'd22
; 
32'd42536: dataIn1 = 32'd23
; 
32'd42537: dataIn1 = 32'd24
; 
32'd42538: dataIn1 = 32'd25
; 
32'd42539: dataIn1 = 32'd27
; 
32'd42540: dataIn1 = 32'd28
; 
32'd42541: dataIn1 = 32'd29
; 
32'd42542: dataIn1 = 32'd30
; 
32'd42543: dataIn1 = 32'd31
; 
32'd42544: dataIn1 = 32'd32
; 
32'd42545: dataIn1 = 32'd33
; 
32'd42546: dataIn1 = 32'd34
; 
32'd42547: dataIn1 = 32'd35
; 
32'd42548: dataIn1 = 32'd37
; 
32'd42549: dataIn1 = 32'd38
; 
32'd42550: dataIn1 = 32'd39
; 
32'd42551: dataIn1 = 32'd40
; 
32'd42552: dataIn1 = 32'd42
; 
32'd42553: dataIn1 = 32'd43
; 
32'd42554: dataIn1 = 32'd44
; 
32'd42555: dataIn1 = 32'd45
; 
32'd42556: dataIn1 = 32'd46
; 
32'd42557: dataIn1 = 32'd47
; 
32'd42558: dataIn1 = 32'd48
; 
32'd42559: dataIn1 = 32'd51
; 
32'd42560: dataIn1 = 32'd52
; 
32'd42561: dataIn1 = 32'd54
; 
32'd42562: dataIn1 = 32'd55
; 
32'd42563: dataIn1 = 32'd56
; 
32'd42564: dataIn1 = 32'd57
; 
32'd42565: dataIn1 = 32'd58
; 
32'd42566: dataIn1 = 32'd60
; 
32'd42567: dataIn1 = 32'd61
; 
32'd42568: dataIn1 = 32'd62
; 
32'd42569: dataIn1 = 32'd63
; 
32'd42570: dataIn1 = 32'd0
; 
32'd42571: dataIn1 = 32'd1
; 
32'd42572: dataIn1 = 32'd3
; 
32'd42573: dataIn1 = 32'd4
; 
32'd42574: dataIn1 = 32'd5
; 
32'd42575: dataIn1 = 32'd6
; 
32'd42576: dataIn1 = 32'd7
; 
32'd42577: dataIn1 = 32'd8
; 
32'd42578: dataIn1 = 32'd9
; 
32'd42579: dataIn1 = 32'd10
; 
32'd42580: dataIn1 = 32'd11
; 
32'd42581: dataIn1 = 32'd12
; 
32'd42582: dataIn1 = 32'd13
; 
32'd42583: dataIn1 = 32'd14
; 
32'd42584: dataIn1 = 32'd16
; 
32'd42585: dataIn1 = 32'd17
; 
32'd42586: dataIn1 = 32'd18
; 
32'd42587: dataIn1 = 32'd20
; 
32'd42588: dataIn1 = 32'd21
; 
32'd42589: dataIn1 = 32'd22
; 
32'd42590: dataIn1 = 32'd23
; 
32'd42591: dataIn1 = 32'd24
; 
32'd42592: dataIn1 = 32'd25
; 
32'd42593: dataIn1 = 32'd27
; 
32'd42594: dataIn1 = 32'd28
; 
32'd42595: dataIn1 = 32'd29
; 
32'd42596: dataIn1 = 32'd30
; 
32'd42597: dataIn1 = 32'd32
; 
32'd42598: dataIn1 = 32'd33
; 
32'd42599: dataIn1 = 32'd34
; 
32'd42600: dataIn1 = 32'd35
; 
32'd42601: dataIn1 = 32'd36
; 
32'd42602: dataIn1 = 32'd37
; 
32'd42603: dataIn1 = 32'd38
; 
32'd42604: dataIn1 = 32'd39
; 
32'd42605: dataIn1 = 32'd40
; 
32'd42606: dataIn1 = 32'd41
; 
32'd42607: dataIn1 = 32'd42
; 
32'd42608: dataIn1 = 32'd43
; 
32'd42609: dataIn1 = 32'd44
; 
32'd42610: dataIn1 = 32'd45
; 
32'd42611: dataIn1 = 32'd46
; 
32'd42612: dataIn1 = 32'd47
; 
32'd42613: dataIn1 = 32'd48
; 
32'd42614: dataIn1 = 32'd49
; 
32'd42615: dataIn1 = 32'd50
; 
32'd42616: dataIn1 = 32'd51
; 
32'd42617: dataIn1 = 32'd52
; 
32'd42618: dataIn1 = 32'd53
; 
32'd42619: dataIn1 = 32'd54
; 
32'd42620: dataIn1 = 32'd57
; 
32'd42621: dataIn1 = 32'd58
; 
32'd42622: dataIn1 = 32'd60
; 
32'd42623: dataIn1 = 32'd61
; 
32'd42624: dataIn1 = 32'd63
; 
32'd42625: dataIn1 = 32'd0
; 
32'd42626: dataIn1 = 32'd1
; 
32'd42627: dataIn1 = 32'd2
; 
32'd42628: dataIn1 = 32'd5
; 
32'd42629: dataIn1 = 32'd7
; 
32'd42630: dataIn1 = 32'd9
; 
32'd42631: dataIn1 = 32'd10
; 
32'd42632: dataIn1 = 32'd11
; 
32'd42633: dataIn1 = 32'd12
; 
32'd42634: dataIn1 = 32'd14
; 
32'd42635: dataIn1 = 32'd15
; 
32'd42636: dataIn1 = 32'd16
; 
32'd42637: dataIn1 = 32'd17
; 
32'd42638: dataIn1 = 32'd18
; 
32'd42639: dataIn1 = 32'd19
; 
32'd42640: dataIn1 = 32'd20
; 
32'd42641: dataIn1 = 32'd21
; 
32'd42642: dataIn1 = 32'd22
; 
32'd42643: dataIn1 = 32'd23
; 
32'd42644: dataIn1 = 32'd24
; 
32'd42645: dataIn1 = 32'd25
; 
32'd42646: dataIn1 = 32'd26
; 
32'd42647: dataIn1 = 32'd27
; 
32'd42648: dataIn1 = 32'd29
; 
32'd42649: dataIn1 = 32'd30
; 
32'd42650: dataIn1 = 32'd31
; 
32'd42651: dataIn1 = 32'd32
; 
32'd42652: dataIn1 = 32'd33
; 
32'd42653: dataIn1 = 32'd34
; 
32'd42654: dataIn1 = 32'd35
; 
32'd42655: dataIn1 = 32'd36
; 
32'd42656: dataIn1 = 32'd37
; 
32'd42657: dataIn1 = 32'd38
; 
32'd42658: dataIn1 = 32'd39
; 
32'd42659: dataIn1 = 32'd40
; 
32'd42660: dataIn1 = 32'd42
; 
32'd42661: dataIn1 = 32'd44
; 
32'd42662: dataIn1 = 32'd45
; 
32'd42663: dataIn1 = 32'd48
; 
32'd42664: dataIn1 = 32'd49
; 
32'd42665: dataIn1 = 32'd50
; 
32'd42666: dataIn1 = 32'd52
; 
32'd42667: dataIn1 = 32'd54
; 
32'd42668: dataIn1 = 32'd55
; 
32'd42669: dataIn1 = 32'd56
; 
32'd42670: dataIn1 = 32'd57
; 
32'd42671: dataIn1 = 32'd58
; 
32'd42672: dataIn1 = 32'd59
; 
32'd42673: dataIn1 = 32'd60
; 
32'd42674: dataIn1 = 32'd61
; 
32'd42675: dataIn1 = 32'd62
; 
32'd42676: dataIn1 = 32'd63
; 
32'd42677: dataIn1 = 32'd0
; 
32'd42678: dataIn1 = 32'd1
; 
32'd42679: dataIn1 = 32'd2
; 
32'd42680: dataIn1 = 32'd3
; 
32'd42681: dataIn1 = 32'd5
; 
32'd42682: dataIn1 = 32'd6
; 
32'd42683: dataIn1 = 32'd7
; 
32'd42684: dataIn1 = 32'd8
; 
32'd42685: dataIn1 = 32'd9
; 
32'd42686: dataIn1 = 32'd10
; 
32'd42687: dataIn1 = 32'd11
; 
32'd42688: dataIn1 = 32'd12
; 
32'd42689: dataIn1 = 32'd13
; 
32'd42690: dataIn1 = 32'd14
; 
32'd42691: dataIn1 = 32'd15
; 
32'd42692: dataIn1 = 32'd16
; 
32'd42693: dataIn1 = 32'd17
; 
32'd42694: dataIn1 = 32'd18
; 
32'd42695: dataIn1 = 32'd19
; 
32'd42696: dataIn1 = 32'd20
; 
32'd42697: dataIn1 = 32'd21
; 
32'd42698: dataIn1 = 32'd22
; 
32'd42699: dataIn1 = 32'd23
; 
32'd42700: dataIn1 = 32'd25
; 
32'd42701: dataIn1 = 32'd26
; 
32'd42702: dataIn1 = 32'd27
; 
32'd42703: dataIn1 = 32'd28
; 
32'd42704: dataIn1 = 32'd29
; 
32'd42705: dataIn1 = 32'd31
; 
32'd42706: dataIn1 = 32'd32
; 
32'd42707: dataIn1 = 32'd33
; 
32'd42708: dataIn1 = 32'd34
; 
32'd42709: dataIn1 = 32'd35
; 
32'd42710: dataIn1 = 32'd36
; 
32'd42711: dataIn1 = 32'd37
; 
32'd42712: dataIn1 = 32'd38
; 
32'd42713: dataIn1 = 32'd39
; 
32'd42714: dataIn1 = 32'd40
; 
32'd42715: dataIn1 = 32'd41
; 
32'd42716: dataIn1 = 32'd42
; 
32'd42717: dataIn1 = 32'd43
; 
32'd42718: dataIn1 = 32'd44
; 
32'd42719: dataIn1 = 32'd45
; 
32'd42720: dataIn1 = 32'd46
; 
32'd42721: dataIn1 = 32'd47
; 
32'd42722: dataIn1 = 32'd48
; 
32'd42723: dataIn1 = 32'd49
; 
32'd42724: dataIn1 = 32'd50
; 
32'd42725: dataIn1 = 32'd51
; 
32'd42726: dataIn1 = 32'd52
; 
32'd42727: dataIn1 = 32'd53
; 
32'd42728: dataIn1 = 32'd55
; 
32'd42729: dataIn1 = 32'd56
; 
32'd42730: dataIn1 = 32'd57
; 
32'd42731: dataIn1 = 32'd58
; 
32'd42732: dataIn1 = 32'd59
; 
32'd42733: dataIn1 = 32'd60
; 
32'd42734: dataIn1 = 32'd61
; 
32'd42735: dataIn1 = 32'd62
; 
32'd42736: dataIn1 = 32'd63
; 
32'd42737: dataIn1 = 32'd0
; 
32'd42738: dataIn1 = 32'd1
; 
32'd42739: dataIn1 = 32'd2
; 
32'd42740: dataIn1 = 32'd5
; 
32'd42741: dataIn1 = 32'd6
; 
32'd42742: dataIn1 = 32'd7
; 
32'd42743: dataIn1 = 32'd9
; 
32'd42744: dataIn1 = 32'd10
; 
32'd42745: dataIn1 = 32'd11
; 
32'd42746: dataIn1 = 32'd13
; 
32'd42747: dataIn1 = 32'd14
; 
32'd42748: dataIn1 = 32'd15
; 
32'd42749: dataIn1 = 32'd16
; 
32'd42750: dataIn1 = 32'd17
; 
32'd42751: dataIn1 = 32'd18
; 
32'd42752: dataIn1 = 32'd19
; 
32'd42753: dataIn1 = 32'd20
; 
32'd42754: dataIn1 = 32'd21
; 
32'd42755: dataIn1 = 32'd22
; 
32'd42756: dataIn1 = 32'd23
; 
32'd42757: dataIn1 = 32'd24
; 
32'd42758: dataIn1 = 32'd25
; 
32'd42759: dataIn1 = 32'd26
; 
32'd42760: dataIn1 = 32'd27
; 
32'd42761: dataIn1 = 32'd28
; 
32'd42762: dataIn1 = 32'd29
; 
32'd42763: dataIn1 = 32'd30
; 
32'd42764: dataIn1 = 32'd31
; 
32'd42765: dataIn1 = 32'd32
; 
32'd42766: dataIn1 = 32'd33
; 
32'd42767: dataIn1 = 32'd34
; 
32'd42768: dataIn1 = 32'd35
; 
32'd42769: dataIn1 = 32'd36
; 
32'd42770: dataIn1 = 32'd37
; 
32'd42771: dataIn1 = 32'd38
; 
32'd42772: dataIn1 = 32'd39
; 
32'd42773: dataIn1 = 32'd40
; 
32'd42774: dataIn1 = 32'd41
; 
32'd42775: dataIn1 = 32'd42
; 
32'd42776: dataIn1 = 32'd43
; 
32'd42777: dataIn1 = 32'd45
; 
32'd42778: dataIn1 = 32'd46
; 
32'd42779: dataIn1 = 32'd47
; 
32'd42780: dataIn1 = 32'd48
; 
32'd42781: dataIn1 = 32'd49
; 
32'd42782: dataIn1 = 32'd50
; 
32'd42783: dataIn1 = 32'd51
; 
32'd42784: dataIn1 = 32'd52
; 
32'd42785: dataIn1 = 32'd53
; 
32'd42786: dataIn1 = 32'd54
; 
32'd42787: dataIn1 = 32'd56
; 
32'd42788: dataIn1 = 32'd57
; 
32'd42789: dataIn1 = 32'd59
; 
32'd42790: dataIn1 = 32'd60
; 
32'd42791: dataIn1 = 32'd61
; 
32'd42792: dataIn1 = 32'd62
; 
32'd42793: dataIn1 = 32'd63
; 
32'd42794: dataIn1 = 32'd0
; 
32'd42795: dataIn1 = 32'd1
; 
32'd42796: dataIn1 = 32'd2
; 
32'd42797: dataIn1 = 32'd3
; 
32'd42798: dataIn1 = 32'd4
; 
32'd42799: dataIn1 = 32'd5
; 
32'd42800: dataIn1 = 32'd6
; 
32'd42801: dataIn1 = 32'd8
; 
32'd42802: dataIn1 = 32'd9
; 
32'd42803: dataIn1 = 32'd10
; 
32'd42804: dataIn1 = 32'd11
; 
32'd42805: dataIn1 = 32'd12
; 
32'd42806: dataIn1 = 32'd14
; 
32'd42807: dataIn1 = 32'd15
; 
32'd42808: dataIn1 = 32'd16
; 
32'd42809: dataIn1 = 32'd17
; 
32'd42810: dataIn1 = 32'd18
; 
32'd42811: dataIn1 = 32'd19
; 
32'd42812: dataIn1 = 32'd20
; 
32'd42813: dataIn1 = 32'd21
; 
32'd42814: dataIn1 = 32'd22
; 
32'd42815: dataIn1 = 32'd23
; 
32'd42816: dataIn1 = 32'd25
; 
32'd42817: dataIn1 = 32'd26
; 
32'd42818: dataIn1 = 32'd27
; 
32'd42819: dataIn1 = 32'd28
; 
32'd42820: dataIn1 = 32'd29
; 
32'd42821: dataIn1 = 32'd31
; 
32'd42822: dataIn1 = 32'd32
; 
32'd42823: dataIn1 = 32'd33
; 
32'd42824: dataIn1 = 32'd34
; 
32'd42825: dataIn1 = 32'd35
; 
32'd42826: dataIn1 = 32'd37
; 
32'd42827: dataIn1 = 32'd39
; 
32'd42828: dataIn1 = 32'd40
; 
32'd42829: dataIn1 = 32'd41
; 
32'd42830: dataIn1 = 32'd42
; 
32'd42831: dataIn1 = 32'd43
; 
32'd42832: dataIn1 = 32'd44
; 
32'd42833: dataIn1 = 32'd45
; 
32'd42834: dataIn1 = 32'd47
; 
32'd42835: dataIn1 = 32'd48
; 
32'd42836: dataIn1 = 32'd50
; 
32'd42837: dataIn1 = 32'd51
; 
32'd42838: dataIn1 = 32'd52
; 
32'd42839: dataIn1 = 32'd53
; 
32'd42840: dataIn1 = 32'd55
; 
32'd42841: dataIn1 = 32'd56
; 
32'd42842: dataIn1 = 32'd57
; 
32'd42843: dataIn1 = 32'd58
; 
32'd42844: dataIn1 = 32'd59
; 
32'd42845: dataIn1 = 32'd60
; 
32'd42846: dataIn1 = 32'd61
; 
32'd42847: dataIn1 = 32'd62
; 
32'd42848: dataIn1 = 32'd63
; 
32'd42849: dataIn1 = 32'd0
; 
32'd42850: dataIn1 = 32'd1
; 
32'd42851: dataIn1 = 32'd2
; 
32'd42852: dataIn1 = 32'd3
; 
32'd42853: dataIn1 = 32'd4
; 
32'd42854: dataIn1 = 32'd5
; 
32'd42855: dataIn1 = 32'd6
; 
32'd42856: dataIn1 = 32'd7
; 
32'd42857: dataIn1 = 32'd10
; 
32'd42858: dataIn1 = 32'd12
; 
32'd42859: dataIn1 = 32'd13
; 
32'd42860: dataIn1 = 32'd15
; 
32'd42861: dataIn1 = 32'd16
; 
32'd42862: dataIn1 = 32'd17
; 
32'd42863: dataIn1 = 32'd18
; 
32'd42864: dataIn1 = 32'd19
; 
32'd42865: dataIn1 = 32'd20
; 
32'd42866: dataIn1 = 32'd22
; 
32'd42867: dataIn1 = 32'd23
; 
32'd42868: dataIn1 = 32'd25
; 
32'd42869: dataIn1 = 32'd26
; 
32'd42870: dataIn1 = 32'd27
; 
32'd42871: dataIn1 = 32'd28
; 
32'd42872: dataIn1 = 32'd29
; 
32'd42873: dataIn1 = 32'd30
; 
32'd42874: dataIn1 = 32'd31
; 
32'd42875: dataIn1 = 32'd32
; 
32'd42876: dataIn1 = 32'd33
; 
32'd42877: dataIn1 = 32'd34
; 
32'd42878: dataIn1 = 32'd35
; 
32'd42879: dataIn1 = 32'd36
; 
32'd42880: dataIn1 = 32'd37
; 
32'd42881: dataIn1 = 32'd38
; 
32'd42882: dataIn1 = 32'd39
; 
32'd42883: dataIn1 = 32'd40
; 
32'd42884: dataIn1 = 32'd41
; 
32'd42885: dataIn1 = 32'd42
; 
32'd42886: dataIn1 = 32'd43
; 
32'd42887: dataIn1 = 32'd44
; 
32'd42888: dataIn1 = 32'd47
; 
32'd42889: dataIn1 = 32'd48
; 
32'd42890: dataIn1 = 32'd49
; 
32'd42891: dataIn1 = 32'd50
; 
32'd42892: dataIn1 = 32'd51
; 
32'd42893: dataIn1 = 32'd52
; 
32'd42894: dataIn1 = 32'd53
; 
32'd42895: dataIn1 = 32'd54
; 
32'd42896: dataIn1 = 32'd55
; 
32'd42897: dataIn1 = 32'd57
; 
32'd42898: dataIn1 = 32'd58
; 
32'd42899: dataIn1 = 32'd59
; 
32'd42900: dataIn1 = 32'd61
; 
32'd42901: dataIn1 = 32'd62
; 
32'd42902: dataIn1 = 32'd63
; 
32'd42903: dataIn1 = 32'd0
; 
32'd42904: dataIn1 = 32'd1
; 
32'd42905: dataIn1 = 32'd2
; 
32'd42906: dataIn1 = 32'd3
; 
32'd42907: dataIn1 = 32'd5
; 
32'd42908: dataIn1 = 32'd6
; 
32'd42909: dataIn1 = 32'd7
; 
32'd42910: dataIn1 = 32'd8
; 
32'd42911: dataIn1 = 32'd9
; 
32'd42912: dataIn1 = 32'd10
; 
32'd42913: dataIn1 = 32'd12
; 
32'd42914: dataIn1 = 32'd14
; 
32'd42915: dataIn1 = 32'd15
; 
32'd42916: dataIn1 = 32'd16
; 
32'd42917: dataIn1 = 32'd18
; 
32'd42918: dataIn1 = 32'd19
; 
32'd42919: dataIn1 = 32'd21
; 
32'd42920: dataIn1 = 32'd22
; 
32'd42921: dataIn1 = 32'd23
; 
32'd42922: dataIn1 = 32'd24
; 
32'd42923: dataIn1 = 32'd25
; 
32'd42924: dataIn1 = 32'd26
; 
32'd42925: dataIn1 = 32'd27
; 
32'd42926: dataIn1 = 32'd28
; 
32'd42927: dataIn1 = 32'd29
; 
32'd42928: dataIn1 = 32'd30
; 
32'd42929: dataIn1 = 32'd31
; 
32'd42930: dataIn1 = 32'd32
; 
32'd42931: dataIn1 = 32'd33
; 
32'd42932: dataIn1 = 32'd34
; 
32'd42933: dataIn1 = 32'd35
; 
32'd42934: dataIn1 = 32'd36
; 
32'd42935: dataIn1 = 32'd37
; 
32'd42936: dataIn1 = 32'd38
; 
32'd42937: dataIn1 = 32'd39
; 
32'd42938: dataIn1 = 32'd40
; 
32'd42939: dataIn1 = 32'd41
; 
32'd42940: dataIn1 = 32'd42
; 
32'd42941: dataIn1 = 32'd43
; 
32'd42942: dataIn1 = 32'd44
; 
32'd42943: dataIn1 = 32'd45
; 
32'd42944: dataIn1 = 32'd46
; 
32'd42945: dataIn1 = 32'd47
; 
32'd42946: dataIn1 = 32'd48
; 
32'd42947: dataIn1 = 32'd49
; 
32'd42948: dataIn1 = 32'd50
; 
32'd42949: dataIn1 = 32'd51
; 
32'd42950: dataIn1 = 32'd52
; 
32'd42951: dataIn1 = 32'd53
; 
32'd42952: dataIn1 = 32'd55
; 
32'd42953: dataIn1 = 32'd56
; 
32'd42954: dataIn1 = 32'd57
; 
32'd42955: dataIn1 = 32'd59
; 
32'd42956: dataIn1 = 32'd60
; 
32'd42957: dataIn1 = 32'd61
; 
32'd42958: dataIn1 = 32'd62
; 
32'd42959: dataIn1 = 32'd0
; 
32'd42960: dataIn1 = 32'd1
; 
32'd42961: dataIn1 = 32'd3
; 
32'd42962: dataIn1 = 32'd4
; 
32'd42963: dataIn1 = 32'd5
; 
32'd42964: dataIn1 = 32'd6
; 
32'd42965: dataIn1 = 32'd7
; 
32'd42966: dataIn1 = 32'd8
; 
32'd42967: dataIn1 = 32'd9
; 
32'd42968: dataIn1 = 32'd10
; 
32'd42969: dataIn1 = 32'd11
; 
32'd42970: dataIn1 = 32'd12
; 
32'd42971: dataIn1 = 32'd13
; 
32'd42972: dataIn1 = 32'd14
; 
32'd42973: dataIn1 = 32'd15
; 
32'd42974: dataIn1 = 32'd17
; 
32'd42975: dataIn1 = 32'd18
; 
32'd42976: dataIn1 = 32'd19
; 
32'd42977: dataIn1 = 32'd20
; 
32'd42978: dataIn1 = 32'd21
; 
32'd42979: dataIn1 = 32'd22
; 
32'd42980: dataIn1 = 32'd23
; 
32'd42981: dataIn1 = 32'd24
; 
32'd42982: dataIn1 = 32'd25
; 
32'd42983: dataIn1 = 32'd26
; 
32'd42984: dataIn1 = 32'd27
; 
32'd42985: dataIn1 = 32'd28
; 
32'd42986: dataIn1 = 32'd29
; 
32'd42987: dataIn1 = 32'd32
; 
32'd42988: dataIn1 = 32'd33
; 
32'd42989: dataIn1 = 32'd34
; 
32'd42990: dataIn1 = 32'd35
; 
32'd42991: dataIn1 = 32'd37
; 
32'd42992: dataIn1 = 32'd38
; 
32'd42993: dataIn1 = 32'd39
; 
32'd42994: dataIn1 = 32'd40
; 
32'd42995: dataIn1 = 32'd41
; 
32'd42996: dataIn1 = 32'd42
; 
32'd42997: dataIn1 = 32'd43
; 
32'd42998: dataIn1 = 32'd44
; 
32'd42999: dataIn1 = 32'd48
; 
32'd43000: dataIn1 = 32'd49
; 
32'd43001: dataIn1 = 32'd50
; 
32'd43002: dataIn1 = 32'd51
; 
32'd43003: dataIn1 = 32'd52
; 
32'd43004: dataIn1 = 32'd53
; 
32'd43005: dataIn1 = 32'd54
; 
32'd43006: dataIn1 = 32'd55
; 
32'd43007: dataIn1 = 32'd56
; 
32'd43008: dataIn1 = 32'd57
; 
32'd43009: dataIn1 = 32'd58
; 
32'd43010: dataIn1 = 32'd59
; 
32'd43011: dataIn1 = 32'd60
; 
32'd43012: dataIn1 = 32'd61
; 
32'd43013: dataIn1 = 32'd62
; 
32'd43014: dataIn1 = 32'd63
; 
32'd43015: dataIn1 = 32'd2
; 
32'd43016: dataIn1 = 32'd4
; 
32'd43017: dataIn1 = 32'd5
; 
32'd43018: dataIn1 = 32'd8
; 
32'd43019: dataIn1 = 32'd9
; 
32'd43020: dataIn1 = 32'd10
; 
32'd43021: dataIn1 = 32'd12
; 
32'd43022: dataIn1 = 32'd15
; 
32'd43023: dataIn1 = 32'd16
; 
32'd43024: dataIn1 = 32'd17
; 
32'd43025: dataIn1 = 32'd18
; 
32'd43026: dataIn1 = 32'd20
; 
32'd43027: dataIn1 = 32'd21
; 
32'd43028: dataIn1 = 32'd22
; 
32'd43029: dataIn1 = 32'd23
; 
32'd43030: dataIn1 = 32'd25
; 
32'd43031: dataIn1 = 32'd28
; 
32'd43032: dataIn1 = 32'd29
; 
32'd43033: dataIn1 = 32'd30
; 
32'd43034: dataIn1 = 32'd31
; 
32'd43035: dataIn1 = 32'd32
; 
32'd43036: dataIn1 = 32'd33
; 
32'd43037: dataIn1 = 32'd34
; 
32'd43038: dataIn1 = 32'd35
; 
32'd43039: dataIn1 = 32'd38
; 
32'd43040: dataIn1 = 32'd40
; 
32'd43041: dataIn1 = 32'd41
; 
32'd43042: dataIn1 = 32'd43
; 
32'd43043: dataIn1 = 32'd44
; 
32'd43044: dataIn1 = 32'd47
; 
32'd43045: dataIn1 = 32'd48
; 
32'd43046: dataIn1 = 32'd49
; 
32'd43047: dataIn1 = 32'd50
; 
32'd43048: dataIn1 = 32'd51
; 
32'd43049: dataIn1 = 32'd52
; 
32'd43050: dataIn1 = 32'd53
; 
32'd43051: dataIn1 = 32'd54
; 
32'd43052: dataIn1 = 32'd55
; 
32'd43053: dataIn1 = 32'd56
; 
32'd43054: dataIn1 = 32'd57
; 
32'd43055: dataIn1 = 32'd58
; 
32'd43056: dataIn1 = 32'd59
; 
32'd43057: dataIn1 = 32'd60
; 
32'd43058: dataIn1 = 32'd62
; 
32'd43059: dataIn1 = 32'd63
; 
32'd43060: dataIn1 = 32'd0
; 
32'd43061: dataIn1 = 32'd1
; 
32'd43062: dataIn1 = 32'd2
; 
32'd43063: dataIn1 = 32'd3
; 
32'd43064: dataIn1 = 32'd4
; 
32'd43065: dataIn1 = 32'd5
; 
32'd43066: dataIn1 = 32'd6
; 
32'd43067: dataIn1 = 32'd7
; 
32'd43068: dataIn1 = 32'd8
; 
32'd43069: dataIn1 = 32'd9
; 
32'd43070: dataIn1 = 32'd10
; 
32'd43071: dataIn1 = 32'd11
; 
32'd43072: dataIn1 = 32'd12
; 
32'd43073: dataIn1 = 32'd13
; 
32'd43074: dataIn1 = 32'd14
; 
32'd43075: dataIn1 = 32'd15
; 
32'd43076: dataIn1 = 32'd17
; 
32'd43077: dataIn1 = 32'd18
; 
32'd43078: dataIn1 = 32'd19
; 
32'd43079: dataIn1 = 32'd20
; 
32'd43080: dataIn1 = 32'd21
; 
32'd43081: dataIn1 = 32'd22
; 
32'd43082: dataIn1 = 32'd23
; 
32'd43083: dataIn1 = 32'd25
; 
32'd43084: dataIn1 = 32'd26
; 
32'd43085: dataIn1 = 32'd27
; 
32'd43086: dataIn1 = 32'd28
; 
32'd43087: dataIn1 = 32'd29
; 
32'd43088: dataIn1 = 32'd30
; 
32'd43089: dataIn1 = 32'd31
; 
32'd43090: dataIn1 = 32'd33
; 
32'd43091: dataIn1 = 32'd34
; 
32'd43092: dataIn1 = 32'd35
; 
32'd43093: dataIn1 = 32'd36
; 
32'd43094: dataIn1 = 32'd37
; 
32'd43095: dataIn1 = 32'd38
; 
32'd43096: dataIn1 = 32'd39
; 
32'd43097: dataIn1 = 32'd40
; 
32'd43098: dataIn1 = 32'd41
; 
32'd43099: dataIn1 = 32'd42
; 
32'd43100: dataIn1 = 32'd43
; 
32'd43101: dataIn1 = 32'd45
; 
32'd43102: dataIn1 = 32'd48
; 
32'd43103: dataIn1 = 32'd49
; 
32'd43104: dataIn1 = 32'd50
; 
32'd43105: dataIn1 = 32'd51
; 
32'd43106: dataIn1 = 32'd52
; 
32'd43107: dataIn1 = 32'd53
; 
32'd43108: dataIn1 = 32'd54
; 
32'd43109: dataIn1 = 32'd55
; 
32'd43110: dataIn1 = 32'd56
; 
32'd43111: dataIn1 = 32'd57
; 
32'd43112: dataIn1 = 32'd58
; 
32'd43113: dataIn1 = 32'd60
; 
32'd43114: dataIn1 = 32'd62
; 
32'd43115: dataIn1 = 32'd63
; 
32'd43116: dataIn1 = 32'd0
; 
32'd43117: dataIn1 = 32'd1
; 
32'd43118: dataIn1 = 32'd2
; 
32'd43119: dataIn1 = 32'd3
; 
32'd43120: dataIn1 = 32'd4
; 
32'd43121: dataIn1 = 32'd5
; 
32'd43122: dataIn1 = 32'd6
; 
32'd43123: dataIn1 = 32'd9
; 
32'd43124: dataIn1 = 32'd10
; 
32'd43125: dataIn1 = 32'd12
; 
32'd43126: dataIn1 = 32'd13
; 
32'd43127: dataIn1 = 32'd14
; 
32'd43128: dataIn1 = 32'd15
; 
32'd43129: dataIn1 = 32'd16
; 
32'd43130: dataIn1 = 32'd17
; 
32'd43131: dataIn1 = 32'd18
; 
32'd43132: dataIn1 = 32'd19
; 
32'd43133: dataIn1 = 32'd20
; 
32'd43134: dataIn1 = 32'd21
; 
32'd43135: dataIn1 = 32'd22
; 
32'd43136: dataIn1 = 32'd23
; 
32'd43137: dataIn1 = 32'd24
; 
32'd43138: dataIn1 = 32'd25
; 
32'd43139: dataIn1 = 32'd26
; 
32'd43140: dataIn1 = 32'd27
; 
32'd43141: dataIn1 = 32'd28
; 
32'd43142: dataIn1 = 32'd29
; 
32'd43143: dataIn1 = 32'd32
; 
32'd43144: dataIn1 = 32'd33
; 
32'd43145: dataIn1 = 32'd34
; 
32'd43146: dataIn1 = 32'd35
; 
32'd43147: dataIn1 = 32'd38
; 
32'd43148: dataIn1 = 32'd40
; 
32'd43149: dataIn1 = 32'd41
; 
32'd43150: dataIn1 = 32'd42
; 
32'd43151: dataIn1 = 32'd43
; 
32'd43152: dataIn1 = 32'd44
; 
32'd43153: dataIn1 = 32'd45
; 
32'd43154: dataIn1 = 32'd46
; 
32'd43155: dataIn1 = 32'd47
; 
32'd43156: dataIn1 = 32'd48
; 
32'd43157: dataIn1 = 32'd49
; 
32'd43158: dataIn1 = 32'd50
; 
32'd43159: dataIn1 = 32'd52
; 
32'd43160: dataIn1 = 32'd53
; 
32'd43161: dataIn1 = 32'd54
; 
32'd43162: dataIn1 = 32'd55
; 
32'd43163: dataIn1 = 32'd56
; 
32'd43164: dataIn1 = 32'd58
; 
32'd43165: dataIn1 = 32'd60
; 
32'd43166: dataIn1 = 32'd61
; 
32'd43167: dataIn1 = 32'd62
; 
32'd43168: dataIn1 = 32'd0
; 
32'd43169: dataIn1 = 32'd1
; 
32'd43170: dataIn1 = 32'd2
; 
32'd43171: dataIn1 = 32'd3
; 
32'd43172: dataIn1 = 32'd5
; 
32'd43173: dataIn1 = 32'd6
; 
32'd43174: dataIn1 = 32'd7
; 
32'd43175: dataIn1 = 32'd8
; 
32'd43176: dataIn1 = 32'd9
; 
32'd43177: dataIn1 = 32'd10
; 
32'd43178: dataIn1 = 32'd11
; 
32'd43179: dataIn1 = 32'd12
; 
32'd43180: dataIn1 = 32'd13
; 
32'd43181: dataIn1 = 32'd14
; 
32'd43182: dataIn1 = 32'd15
; 
32'd43183: dataIn1 = 32'd16
; 
32'd43184: dataIn1 = 32'd17
; 
32'd43185: dataIn1 = 32'd18
; 
32'd43186: dataIn1 = 32'd20
; 
32'd43187: dataIn1 = 32'd21
; 
32'd43188: dataIn1 = 32'd22
; 
32'd43189: dataIn1 = 32'd23
; 
32'd43190: dataIn1 = 32'd24
; 
32'd43191: dataIn1 = 32'd25
; 
32'd43192: dataIn1 = 32'd26
; 
32'd43193: dataIn1 = 32'd27
; 
32'd43194: dataIn1 = 32'd28
; 
32'd43195: dataIn1 = 32'd29
; 
32'd43196: dataIn1 = 32'd30
; 
32'd43197: dataIn1 = 32'd31
; 
32'd43198: dataIn1 = 32'd32
; 
32'd43199: dataIn1 = 32'd33
; 
32'd43200: dataIn1 = 32'd34
; 
32'd43201: dataIn1 = 32'd35
; 
32'd43202: dataIn1 = 32'd36
; 
32'd43203: dataIn1 = 32'd37
; 
32'd43204: dataIn1 = 32'd39
; 
32'd43205: dataIn1 = 32'd40
; 
32'd43206: dataIn1 = 32'd41
; 
32'd43207: dataIn1 = 32'd42
; 
32'd43208: dataIn1 = 32'd43
; 
32'd43209: dataIn1 = 32'd44
; 
32'd43210: dataIn1 = 32'd45
; 
32'd43211: dataIn1 = 32'd46
; 
32'd43212: dataIn1 = 32'd47
; 
32'd43213: dataIn1 = 32'd48
; 
32'd43214: dataIn1 = 32'd49
; 
32'd43215: dataIn1 = 32'd51
; 
32'd43216: dataIn1 = 32'd52
; 
32'd43217: dataIn1 = 32'd53
; 
32'd43218: dataIn1 = 32'd54
; 
32'd43219: dataIn1 = 32'd55
; 
32'd43220: dataIn1 = 32'd56
; 
32'd43221: dataIn1 = 32'd57
; 
32'd43222: dataIn1 = 32'd58
; 
32'd43223: dataIn1 = 32'd59
; 
32'd43224: dataIn1 = 32'd60
; 
32'd43225: dataIn1 = 32'd62
; 
32'd43226: dataIn1 = 32'd0
; 
32'd43227: dataIn1 = 32'd1
; 
32'd43228: dataIn1 = 32'd2
; 
32'd43229: dataIn1 = 32'd4
; 
32'd43230: dataIn1 = 32'd5
; 
32'd43231: dataIn1 = 32'd6
; 
32'd43232: dataIn1 = 32'd7
; 
32'd43233: dataIn1 = 32'd8
; 
32'd43234: dataIn1 = 32'd9
; 
32'd43235: dataIn1 = 32'd10
; 
32'd43236: dataIn1 = 32'd11
; 
32'd43237: dataIn1 = 32'd12
; 
32'd43238: dataIn1 = 32'd13
; 
32'd43239: dataIn1 = 32'd14
; 
32'd43240: dataIn1 = 32'd15
; 
32'd43241: dataIn1 = 32'd16
; 
32'd43242: dataIn1 = 32'd17
; 
32'd43243: dataIn1 = 32'd18
; 
32'd43244: dataIn1 = 32'd20
; 
32'd43245: dataIn1 = 32'd21
; 
32'd43246: dataIn1 = 32'd22
; 
32'd43247: dataIn1 = 32'd23
; 
32'd43248: dataIn1 = 32'd24
; 
32'd43249: dataIn1 = 32'd25
; 
32'd43250: dataIn1 = 32'd26
; 
32'd43251: dataIn1 = 32'd27
; 
32'd43252: dataIn1 = 32'd28
; 
32'd43253: dataIn1 = 32'd29
; 
32'd43254: dataIn1 = 32'd30
; 
32'd43255: dataIn1 = 32'd31
; 
32'd43256: dataIn1 = 32'd32
; 
32'd43257: dataIn1 = 32'd33
; 
32'd43258: dataIn1 = 32'd34
; 
32'd43259: dataIn1 = 32'd35
; 
32'd43260: dataIn1 = 32'd36
; 
32'd43261: dataIn1 = 32'd37
; 
32'd43262: dataIn1 = 32'd38
; 
32'd43263: dataIn1 = 32'd39
; 
32'd43264: dataIn1 = 32'd40
; 
32'd43265: dataIn1 = 32'd41
; 
32'd43266: dataIn1 = 32'd42
; 
32'd43267: dataIn1 = 32'd43
; 
32'd43268: dataIn1 = 32'd44
; 
32'd43269: dataIn1 = 32'd45
; 
32'd43270: dataIn1 = 32'd46
; 
32'd43271: dataIn1 = 32'd47
; 
32'd43272: dataIn1 = 32'd48
; 
32'd43273: dataIn1 = 32'd49
; 
32'd43274: dataIn1 = 32'd50
; 
32'd43275: dataIn1 = 32'd52
; 
32'd43276: dataIn1 = 32'd53
; 
32'd43277: dataIn1 = 32'd54
; 
32'd43278: dataIn1 = 32'd55
; 
32'd43279: dataIn1 = 32'd56
; 
32'd43280: dataIn1 = 32'd57
; 
32'd43281: dataIn1 = 32'd59
; 
32'd43282: dataIn1 = 32'd60
; 
32'd43283: dataIn1 = 32'd61
; 
32'd43284: dataIn1 = 32'd0
; 
32'd43285: dataIn1 = 32'd1
; 
32'd43286: dataIn1 = 32'd3
; 
32'd43287: dataIn1 = 32'd4
; 
32'd43288: dataIn1 = 32'd5
; 
32'd43289: dataIn1 = 32'd6
; 
32'd43290: dataIn1 = 32'd7
; 
32'd43291: dataIn1 = 32'd8
; 
32'd43292: dataIn1 = 32'd9
; 
32'd43293: dataIn1 = 32'd10
; 
32'd43294: dataIn1 = 32'd11
; 
32'd43295: dataIn1 = 32'd12
; 
32'd43296: dataIn1 = 32'd13
; 
32'd43297: dataIn1 = 32'd14
; 
32'd43298: dataIn1 = 32'd15
; 
32'd43299: dataIn1 = 32'd16
; 
32'd43300: dataIn1 = 32'd17
; 
32'd43301: dataIn1 = 32'd18
; 
32'd43302: dataIn1 = 32'd19
; 
32'd43303: dataIn1 = 32'd20
; 
32'd43304: dataIn1 = 32'd22
; 
32'd43305: dataIn1 = 32'd23
; 
32'd43306: dataIn1 = 32'd25
; 
32'd43307: dataIn1 = 32'd26
; 
32'd43308: dataIn1 = 32'd29
; 
32'd43309: dataIn1 = 32'd30
; 
32'd43310: dataIn1 = 32'd33
; 
32'd43311: dataIn1 = 32'd34
; 
32'd43312: dataIn1 = 32'd35
; 
32'd43313: dataIn1 = 32'd36
; 
32'd43314: dataIn1 = 32'd37
; 
32'd43315: dataIn1 = 32'd38
; 
32'd43316: dataIn1 = 32'd41
; 
32'd43317: dataIn1 = 32'd42
; 
32'd43318: dataIn1 = 32'd44
; 
32'd43319: dataIn1 = 32'd45
; 
32'd43320: dataIn1 = 32'd46
; 
32'd43321: dataIn1 = 32'd48
; 
32'd43322: dataIn1 = 32'd49
; 
32'd43323: dataIn1 = 32'd51
; 
32'd43324: dataIn1 = 32'd52
; 
32'd43325: dataIn1 = 32'd54
; 
32'd43326: dataIn1 = 32'd55
; 
32'd43327: dataIn1 = 32'd57
; 
32'd43328: dataIn1 = 32'd58
; 
32'd43329: dataIn1 = 32'd59
; 
32'd43330: dataIn1 = 32'd60
; 
32'd43331: dataIn1 = 32'd61
; 
32'd43332: dataIn1 = 32'd62
; 
32'd43333: dataIn1 = 32'd63
; 
32'd43334: dataIn1 = 32'd0
; 
32'd43335: dataIn1 = 32'd3
; 
32'd43336: dataIn1 = 32'd4
; 
32'd43337: dataIn1 = 32'd5
; 
32'd43338: dataIn1 = 32'd6
; 
32'd43339: dataIn1 = 32'd7
; 
32'd43340: dataIn1 = 32'd8
; 
32'd43341: dataIn1 = 32'd9
; 
32'd43342: dataIn1 = 32'd10
; 
32'd43343: dataIn1 = 32'd11
; 
32'd43344: dataIn1 = 32'd12
; 
32'd43345: dataIn1 = 32'd13
; 
32'd43346: dataIn1 = 32'd14
; 
32'd43347: dataIn1 = 32'd15
; 
32'd43348: dataIn1 = 32'd16
; 
32'd43349: dataIn1 = 32'd17
; 
32'd43350: dataIn1 = 32'd18
; 
32'd43351: dataIn1 = 32'd19
; 
32'd43352: dataIn1 = 32'd20
; 
32'd43353: dataIn1 = 32'd21
; 
32'd43354: dataIn1 = 32'd22
; 
32'd43355: dataIn1 = 32'd23
; 
32'd43356: dataIn1 = 32'd25
; 
32'd43357: dataIn1 = 32'd26
; 
32'd43358: dataIn1 = 32'd27
; 
32'd43359: dataIn1 = 32'd28
; 
32'd43360: dataIn1 = 32'd29
; 
32'd43361: dataIn1 = 32'd30
; 
32'd43362: dataIn1 = 32'd31
; 
32'd43363: dataIn1 = 32'd32
; 
32'd43364: dataIn1 = 32'd33
; 
32'd43365: dataIn1 = 32'd34
; 
32'd43366: dataIn1 = 32'd35
; 
32'd43367: dataIn1 = 32'd36
; 
32'd43368: dataIn1 = 32'd37
; 
32'd43369: dataIn1 = 32'd38
; 
32'd43370: dataIn1 = 32'd39
; 
32'd43371: dataIn1 = 32'd40
; 
32'd43372: dataIn1 = 32'd42
; 
32'd43373: dataIn1 = 32'd43
; 
32'd43374: dataIn1 = 32'd46
; 
32'd43375: dataIn1 = 32'd47
; 
32'd43376: dataIn1 = 32'd48
; 
32'd43377: dataIn1 = 32'd49
; 
32'd43378: dataIn1 = 32'd50
; 
32'd43379: dataIn1 = 32'd51
; 
32'd43380: dataIn1 = 32'd52
; 
32'd43381: dataIn1 = 32'd53
; 
32'd43382: dataIn1 = 32'd54
; 
32'd43383: dataIn1 = 32'd55
; 
32'd43384: dataIn1 = 32'd56
; 
32'd43385: dataIn1 = 32'd58
; 
32'd43386: dataIn1 = 32'd59
; 
32'd43387: dataIn1 = 32'd60
; 
32'd43388: dataIn1 = 32'd61
; 
32'd43389: dataIn1 = 32'd62
; 
32'd43390: dataIn1 = 32'd63
; 
32'd43391: dataIn1 = 32'd0
; 
32'd43392: dataIn1 = 32'd1
; 
32'd43393: dataIn1 = 32'd2
; 
32'd43394: dataIn1 = 32'd3
; 
32'd43395: dataIn1 = 32'd4
; 
32'd43396: dataIn1 = 32'd5
; 
32'd43397: dataIn1 = 32'd6
; 
32'd43398: dataIn1 = 32'd7
; 
32'd43399: dataIn1 = 32'd8
; 
32'd43400: dataIn1 = 32'd9
; 
32'd43401: dataIn1 = 32'd11
; 
32'd43402: dataIn1 = 32'd13
; 
32'd43403: dataIn1 = 32'd14
; 
32'd43404: dataIn1 = 32'd15
; 
32'd43405: dataIn1 = 32'd16
; 
32'd43406: dataIn1 = 32'd17
; 
32'd43407: dataIn1 = 32'd19
; 
32'd43408: dataIn1 = 32'd20
; 
32'd43409: dataIn1 = 32'd23
; 
32'd43410: dataIn1 = 32'd24
; 
32'd43411: dataIn1 = 32'd25
; 
32'd43412: dataIn1 = 32'd26
; 
32'd43413: dataIn1 = 32'd27
; 
32'd43414: dataIn1 = 32'd28
; 
32'd43415: dataIn1 = 32'd29
; 
32'd43416: dataIn1 = 32'd30
; 
32'd43417: dataIn1 = 32'd31
; 
32'd43418: dataIn1 = 32'd32
; 
32'd43419: dataIn1 = 32'd33
; 
32'd43420: dataIn1 = 32'd34
; 
32'd43421: dataIn1 = 32'd35
; 
32'd43422: dataIn1 = 32'd36
; 
32'd43423: dataIn1 = 32'd37
; 
32'd43424: dataIn1 = 32'd38
; 
32'd43425: dataIn1 = 32'd40
; 
32'd43426: dataIn1 = 32'd41
; 
32'd43427: dataIn1 = 32'd42
; 
32'd43428: dataIn1 = 32'd43
; 
32'd43429: dataIn1 = 32'd44
; 
32'd43430: dataIn1 = 32'd45
; 
32'd43431: dataIn1 = 32'd46
; 
32'd43432: dataIn1 = 32'd47
; 
32'd43433: dataIn1 = 32'd49
; 
32'd43434: dataIn1 = 32'd51
; 
32'd43435: dataIn1 = 32'd52
; 
32'd43436: dataIn1 = 32'd53
; 
32'd43437: dataIn1 = 32'd54
; 
32'd43438: dataIn1 = 32'd55
; 
32'd43439: dataIn1 = 32'd56
; 
32'd43440: dataIn1 = 32'd57
; 
32'd43441: dataIn1 = 32'd58
; 
32'd43442: dataIn1 = 32'd59
; 
32'd43443: dataIn1 = 32'd60
; 
32'd43444: dataIn1 = 32'd61
; 
32'd43445: dataIn1 = 32'd62
; 
32'd43446: dataIn1 = 32'd63
; 
32'd43447: dataIn1 = 32'd0
; 
32'd43448: dataIn1 = 32'd1
; 
32'd43449: dataIn1 = 32'd2
; 
32'd43450: dataIn1 = 32'd3
; 
32'd43451: dataIn1 = 32'd4
; 
32'd43452: dataIn1 = 32'd5
; 
32'd43453: dataIn1 = 32'd6
; 
32'd43454: dataIn1 = 32'd7
; 
32'd43455: dataIn1 = 32'd8
; 
32'd43456: dataIn1 = 32'd9
; 
32'd43457: dataIn1 = 32'd10
; 
32'd43458: dataIn1 = 32'd11
; 
32'd43459: dataIn1 = 32'd12
; 
32'd43460: dataIn1 = 32'd13
; 
32'd43461: dataIn1 = 32'd15
; 
32'd43462: dataIn1 = 32'd16
; 
32'd43463: dataIn1 = 32'd17
; 
32'd43464: dataIn1 = 32'd18
; 
32'd43465: dataIn1 = 32'd19
; 
32'd43466: dataIn1 = 32'd20
; 
32'd43467: dataIn1 = 32'd21
; 
32'd43468: dataIn1 = 32'd22
; 
32'd43469: dataIn1 = 32'd25
; 
32'd43470: dataIn1 = 32'd26
; 
32'd43471: dataIn1 = 32'd27
; 
32'd43472: dataIn1 = 32'd28
; 
32'd43473: dataIn1 = 32'd29
; 
32'd43474: dataIn1 = 32'd30
; 
32'd43475: dataIn1 = 32'd31
; 
32'd43476: dataIn1 = 32'd32
; 
32'd43477: dataIn1 = 32'd33
; 
32'd43478: dataIn1 = 32'd34
; 
32'd43479: dataIn1 = 32'd35
; 
32'd43480: dataIn1 = 32'd36
; 
32'd43481: dataIn1 = 32'd37
; 
32'd43482: dataIn1 = 32'd38
; 
32'd43483: dataIn1 = 32'd40
; 
32'd43484: dataIn1 = 32'd41
; 
32'd43485: dataIn1 = 32'd42
; 
32'd43486: dataIn1 = 32'd43
; 
32'd43487: dataIn1 = 32'd45
; 
32'd43488: dataIn1 = 32'd46
; 
32'd43489: dataIn1 = 32'd47
; 
32'd43490: dataIn1 = 32'd48
; 
32'd43491: dataIn1 = 32'd49
; 
32'd43492: dataIn1 = 32'd51
; 
32'd43493: dataIn1 = 32'd52
; 
32'd43494: dataIn1 = 32'd53
; 
32'd43495: dataIn1 = 32'd54
; 
32'd43496: dataIn1 = 32'd55
; 
32'd43497: dataIn1 = 32'd56
; 
32'd43498: dataIn1 = 32'd57
; 
32'd43499: dataIn1 = 32'd58
; 
32'd43500: dataIn1 = 32'd59
; 
32'd43501: dataIn1 = 32'd60
; 
32'd43502: dataIn1 = 32'd61
; 
32'd43503: dataIn1 = 32'd63
; 
32'd43504: dataIn1 = 32'd0
; 
32'd43505: dataIn1 = 32'd1
; 
32'd43506: dataIn1 = 32'd3
; 
32'd43507: dataIn1 = 32'd4
; 
32'd43508: dataIn1 = 32'd5
; 
32'd43509: dataIn1 = 32'd6
; 
32'd43510: dataIn1 = 32'd7
; 
32'd43511: dataIn1 = 32'd8
; 
32'd43512: dataIn1 = 32'd9
; 
32'd43513: dataIn1 = 32'd11
; 
32'd43514: dataIn1 = 32'd12
; 
32'd43515: dataIn1 = 32'd13
; 
32'd43516: dataIn1 = 32'd14
; 
32'd43517: dataIn1 = 32'd15
; 
32'd43518: dataIn1 = 32'd16
; 
32'd43519: dataIn1 = 32'd17
; 
32'd43520: dataIn1 = 32'd19
; 
32'd43521: dataIn1 = 32'd20
; 
32'd43522: dataIn1 = 32'd21
; 
32'd43523: dataIn1 = 32'd22
; 
32'd43524: dataIn1 = 32'd23
; 
32'd43525: dataIn1 = 32'd24
; 
32'd43526: dataIn1 = 32'd25
; 
32'd43527: dataIn1 = 32'd26
; 
32'd43528: dataIn1 = 32'd27
; 
32'd43529: dataIn1 = 32'd28
; 
32'd43530: dataIn1 = 32'd29
; 
32'd43531: dataIn1 = 32'd30
; 
32'd43532: dataIn1 = 32'd31
; 
32'd43533: dataIn1 = 32'd32
; 
32'd43534: dataIn1 = 32'd33
; 
32'd43535: dataIn1 = 32'd34
; 
32'd43536: dataIn1 = 32'd35
; 
32'd43537: dataIn1 = 32'd36
; 
32'd43538: dataIn1 = 32'd37
; 
32'd43539: dataIn1 = 32'd38
; 
32'd43540: dataIn1 = 32'd39
; 
32'd43541: dataIn1 = 32'd40
; 
32'd43542: dataIn1 = 32'd41
; 
32'd43543: dataIn1 = 32'd42
; 
32'd43544: dataIn1 = 32'd43
; 
32'd43545: dataIn1 = 32'd44
; 
32'd43546: dataIn1 = 32'd45
; 
32'd43547: dataIn1 = 32'd46
; 
32'd43548: dataIn1 = 32'd48
; 
32'd43549: dataIn1 = 32'd49
; 
32'd43550: dataIn1 = 32'd50
; 
32'd43551: dataIn1 = 32'd51
; 
32'd43552: dataIn1 = 32'd52
; 
32'd43553: dataIn1 = 32'd53
; 
32'd43554: dataIn1 = 32'd54
; 
32'd43555: dataIn1 = 32'd55
; 
32'd43556: dataIn1 = 32'd57
; 
32'd43557: dataIn1 = 32'd58
; 
32'd43558: dataIn1 = 32'd59
; 
32'd43559: dataIn1 = 32'd60
; 
32'd43560: dataIn1 = 32'd61
; 
32'd43561: dataIn1 = 32'd62
; 
32'd43562: dataIn1 = 32'd63
; 
32'd43563: dataIn1 = 32'd0
; 
32'd43564: dataIn1 = 32'd1
; 
32'd43565: dataIn1 = 32'd2
; 
32'd43566: dataIn1 = 32'd3
; 
32'd43567: dataIn1 = 32'd4
; 
32'd43568: dataIn1 = 32'd5
; 
32'd43569: dataIn1 = 32'd6
; 
32'd43570: dataIn1 = 32'd7
; 
32'd43571: dataIn1 = 32'd8
; 
32'd43572: dataIn1 = 32'd9
; 
32'd43573: dataIn1 = 32'd10
; 
32'd43574: dataIn1 = 32'd11
; 
32'd43575: dataIn1 = 32'd12
; 
32'd43576: dataIn1 = 32'd13
; 
32'd43577: dataIn1 = 32'd14
; 
32'd43578: dataIn1 = 32'd15
; 
32'd43579: dataIn1 = 32'd16
; 
32'd43580: dataIn1 = 32'd17
; 
32'd43581: dataIn1 = 32'd18
; 
32'd43582: dataIn1 = 32'd19
; 
32'd43583: dataIn1 = 32'd20
; 
32'd43584: dataIn1 = 32'd21
; 
32'd43585: dataIn1 = 32'd22
; 
32'd43586: dataIn1 = 32'd23
; 
32'd43587: dataIn1 = 32'd24
; 
32'd43588: dataIn1 = 32'd25
; 
32'd43589: dataIn1 = 32'd26
; 
32'd43590: dataIn1 = 32'd27
; 
32'd43591: dataIn1 = 32'd28
; 
32'd43592: dataIn1 = 32'd29
; 
32'd43593: dataIn1 = 32'd30
; 
32'd43594: dataIn1 = 32'd31
; 
32'd43595: dataIn1 = 32'd32
; 
32'd43596: dataIn1 = 32'd33
; 
32'd43597: dataIn1 = 32'd34
; 
32'd43598: dataIn1 = 32'd35
; 
32'd43599: dataIn1 = 32'd36
; 
32'd43600: dataIn1 = 32'd37
; 
32'd43601: dataIn1 = 32'd39
; 
32'd43602: dataIn1 = 32'd40
; 
32'd43603: dataIn1 = 32'd41
; 
32'd43604: dataIn1 = 32'd42
; 
32'd43605: dataIn1 = 32'd43
; 
32'd43606: dataIn1 = 32'd44
; 
32'd43607: dataIn1 = 32'd45
; 
32'd43608: dataIn1 = 32'd46
; 
32'd43609: dataIn1 = 32'd47
; 
32'd43610: dataIn1 = 32'd48
; 
32'd43611: dataIn1 = 32'd49
; 
32'd43612: dataIn1 = 32'd50
; 
32'd43613: dataIn1 = 32'd51
; 
32'd43614: dataIn1 = 32'd54
; 
32'd43615: dataIn1 = 32'd55
; 
32'd43616: dataIn1 = 32'd56
; 
32'd43617: dataIn1 = 32'd57
; 
32'd43618: dataIn1 = 32'd58
; 
32'd43619: dataIn1 = 32'd59
; 
32'd43620: dataIn1 = 32'd60
; 
32'd43621: dataIn1 = 32'd61
; 
32'd43622: dataIn1 = 32'd62
; 
32'd43623: dataIn1 = 32'd63
; 
32'd43624: dataIn1 = 32'd0
; 
32'd43625: dataIn1 = 32'd2
; 
32'd43626: dataIn1 = 32'd3
; 
32'd43627: dataIn1 = 32'd5
; 
32'd43628: dataIn1 = 32'd7
; 
32'd43629: dataIn1 = 32'd8
; 
32'd43630: dataIn1 = 32'd9
; 
32'd43631: dataIn1 = 32'd10
; 
32'd43632: dataIn1 = 32'd11
; 
32'd43633: dataIn1 = 32'd13
; 
32'd43634: dataIn1 = 32'd14
; 
32'd43635: dataIn1 = 32'd15
; 
32'd43636: dataIn1 = 32'd17
; 
32'd43637: dataIn1 = 32'd18
; 
32'd43638: dataIn1 = 32'd19
; 
32'd43639: dataIn1 = 32'd20
; 
32'd43640: dataIn1 = 32'd22
; 
32'd43641: dataIn1 = 32'd23
; 
32'd43642: dataIn1 = 32'd26
; 
32'd43643: dataIn1 = 32'd28
; 
32'd43644: dataIn1 = 32'd29
; 
32'd43645: dataIn1 = 32'd30
; 
32'd43646: dataIn1 = 32'd31
; 
32'd43647: dataIn1 = 32'd32
; 
32'd43648: dataIn1 = 32'd33
; 
32'd43649: dataIn1 = 32'd34
; 
32'd43650: dataIn1 = 32'd35
; 
32'd43651: dataIn1 = 32'd36
; 
32'd43652: dataIn1 = 32'd37
; 
32'd43653: dataIn1 = 32'd38
; 
32'd43654: dataIn1 = 32'd39
; 
32'd43655: dataIn1 = 32'd40
; 
32'd43656: dataIn1 = 32'd42
; 
32'd43657: dataIn1 = 32'd43
; 
32'd43658: dataIn1 = 32'd44
; 
32'd43659: dataIn1 = 32'd45
; 
32'd43660: dataIn1 = 32'd46
; 
32'd43661: dataIn1 = 32'd47
; 
32'd43662: dataIn1 = 32'd48
; 
32'd43663: dataIn1 = 32'd50
; 
32'd43664: dataIn1 = 32'd51
; 
32'd43665: dataIn1 = 32'd52
; 
32'd43666: dataIn1 = 32'd53
; 
32'd43667: dataIn1 = 32'd54
; 
32'd43668: dataIn1 = 32'd55
; 
32'd43669: dataIn1 = 32'd56
; 
32'd43670: dataIn1 = 32'd57
; 
32'd43671: dataIn1 = 32'd58
; 
32'd43672: dataIn1 = 32'd59
; 
32'd43673: dataIn1 = 32'd60
; 
32'd43674: dataIn1 = 32'd61
; 
32'd43675: dataIn1 = 32'd62
; 
32'd43676: dataIn1 = 32'd0
; 
32'd43677: dataIn1 = 32'd1
; 
32'd43678: dataIn1 = 32'd2
; 
32'd43679: dataIn1 = 32'd3
; 
32'd43680: dataIn1 = 32'd4
; 
32'd43681: dataIn1 = 32'd5
; 
32'd43682: dataIn1 = 32'd6
; 
32'd43683: dataIn1 = 32'd7
; 
32'd43684: dataIn1 = 32'd8
; 
32'd43685: dataIn1 = 32'd9
; 
32'd43686: dataIn1 = 32'd10
; 
32'd43687: dataIn1 = 32'd12
; 
32'd43688: dataIn1 = 32'd13
; 
32'd43689: dataIn1 = 32'd14
; 
32'd43690: dataIn1 = 32'd15
; 
32'd43691: dataIn1 = 32'd16
; 
32'd43692: dataIn1 = 32'd17
; 
32'd43693: dataIn1 = 32'd19
; 
32'd43694: dataIn1 = 32'd20
; 
32'd43695: dataIn1 = 32'd21
; 
32'd43696: dataIn1 = 32'd22
; 
32'd43697: dataIn1 = 32'd23
; 
32'd43698: dataIn1 = 32'd24
; 
32'd43699: dataIn1 = 32'd25
; 
32'd43700: dataIn1 = 32'd27
; 
32'd43701: dataIn1 = 32'd29
; 
32'd43702: dataIn1 = 32'd30
; 
32'd43703: dataIn1 = 32'd32
; 
32'd43704: dataIn1 = 32'd33
; 
32'd43705: dataIn1 = 32'd34
; 
32'd43706: dataIn1 = 32'd35
; 
32'd43707: dataIn1 = 32'd37
; 
32'd43708: dataIn1 = 32'd38
; 
32'd43709: dataIn1 = 32'd39
; 
32'd43710: dataIn1 = 32'd40
; 
32'd43711: dataIn1 = 32'd41
; 
32'd43712: dataIn1 = 32'd42
; 
32'd43713: dataIn1 = 32'd43
; 
32'd43714: dataIn1 = 32'd44
; 
32'd43715: dataIn1 = 32'd45
; 
32'd43716: dataIn1 = 32'd47
; 
32'd43717: dataIn1 = 32'd48
; 
32'd43718: dataIn1 = 32'd49
; 
32'd43719: dataIn1 = 32'd50
; 
32'd43720: dataIn1 = 32'd51
; 
32'd43721: dataIn1 = 32'd52
; 
32'd43722: dataIn1 = 32'd54
; 
32'd43723: dataIn1 = 32'd55
; 
32'd43724: dataIn1 = 32'd56
; 
32'd43725: dataIn1 = 32'd57
; 
32'd43726: dataIn1 = 32'd58
; 
32'd43727: dataIn1 = 32'd59
; 
32'd43728: dataIn1 = 32'd60
; 
32'd43729: dataIn1 = 32'd61
; 
32'd43730: dataIn1 = 32'd63
; 
32'd43731: dataIn1 = 32'd; 
32'd43732: dataIn1 = 32'd; 
32'd43733: dataIn1 = 32'd; 
32'd43734: dataIn1 = 32'd; 
32'd43735: dataIn1 = 32'd; 
32'd43736: dataIn1 = 32'd; 
32'd43737: dataIn1 = 32'd; 
32'd43738: dataIn1 = 32'd; 
32'd43739: dataIn1 = 32'd; 
32'd43740: dataIn1 = 32'd; 
32'd43741: dataIn1 = 32'd; 
32'd43742: dataIn1 = 32'd; 
32'd43743: dataIn1 = 32'd; 
32'd43744: dataIn1 = 32'd; 
32'd43745: dataIn1 = 32'd; 
32'd43746: dataIn1 = 32'd; 
32'd43747: dataIn1 = 32'd; 
32'd43748: dataIn1 = 32'd; 
32'd43749: dataIn1 = 32'd; 
32'd43750: dataIn1 = 32'd; 
32'd43751: dataIn1 = 32'd; 
32'd43752: dataIn1 = 32'd; 
32'd43753: dataIn1 = 32'd; 
32'd43754: dataIn1 = 32'd; 
32'd43755: dataIn1 = 32'd; 
32'd43756: dataIn1 = 32'd; 
32'd43757: dataIn1 = 32'd; 
32'd43758: dataIn1 = 32'd; 
32'd43759: dataIn1 = 32'd; 
32'd43760: dataIn1 = 32'd; 
32'd43761: dataIn1 = 32'd; 
32'd43762: dataIn1 = 32'd; 
32'd43763: dataIn1 = 32'd; 
32'd43764: dataIn1 = 32'd; 
32'd43765: dataIn1 = 32'd; 
32'd43766: dataIn1 = 32'd; 
32'd43767: dataIn1 = 32'd; 
32'd43768: dataIn1 = 32'd; 
32'd43769: dataIn1 = 32'd; 
32'd43770: dataIn1 = 32'd; 
32'd43771: dataIn1 = 32'd; 
32'd43772: dataIn1 = 32'd; 
32'd43773: dataIn1 = 32'd; 
32'd43774: dataIn1 = 32'd; 
32'd43775: dataIn1 = 32'd; 
32'd43776: dataIn1 = 32'd; 
32'd43777: dataIn1 = 32'd; 
32'd43778: dataIn1 = 32'd; 
32'd43779: dataIn1 = 32'd; 
32'd43780: dataIn1 = 32'd; 
32'd43781: dataIn1 = 32'd; 
32'd43782: dataIn1 = 32'd; 
32'd43783: dataIn1 = 32'd; 
32'd43784: dataIn1 = 32'd; 
32'd43785: dataIn1 = 32'd; 
32'd43786: dataIn1 = 32'd; 
32'd43787: dataIn1 = 32'd; 
32'd43788: dataIn1 = 32'd; 
32'd43789: dataIn1 = 32'd; 
32'd43790: dataIn1 = 32'd; 
32'd43791: dataIn1 = 32'd; 
32'd43792: dataIn1 = 32'd; 
32'd43793: dataIn1 = 32'd; 
32'd43794: dataIn1 = 32'd; 
32'd43795: dataIn1 = 32'd; 
32'd43796: dataIn1 = 32'd; 
32'd43797: dataIn1 = 32'd; 
32'd43798: dataIn1 = 32'd; 
32'd43799: dataIn1 = 32'd; 
32'd43800: dataIn1 = 32'd; 
32'd43801: dataIn1 = 32'd; 
32'd43802: dataIn1 = 32'd; 
32'd43803: dataIn1 = 32'd; 
32'd43804: dataIn1 = 32'd; 
32'd43805: dataIn1 = 32'd; 
32'd43806: dataIn1 = 32'd; 
32'd43807: dataIn1 = 32'd; 
32'd43808: dataIn1 = 32'd; 
32'd43809: dataIn1 = 32'd; 
32'd43810: dataIn1 = 32'd; 
32'd43811: dataIn1 = 32'd; 
32'd43812: dataIn1 = 32'd; 
32'd43813: dataIn1 = 32'd; 
32'd43814: dataIn1 = 32'd; 
32'd43815: dataIn1 = 32'd; 
32'd43816: dataIn1 = 32'd; 
32'd43817: dataIn1 = 32'd; 
32'd43818: dataIn1 = 32'd; 
32'd43819: dataIn1 = 32'd; 
32'd43820: dataIn1 = 32'd; 
32'd43821: dataIn1 = 32'd; 
32'd43822: dataIn1 = 32'd; 
32'd43823: dataIn1 = 32'd; 
32'd43824: dataIn1 = 32'd; 
32'd43825: dataIn1 = 32'd; 
32'd43826: dataIn1 = 32'd; 
32'd43827: dataIn1 = 32'd; 
32'd43828: dataIn1 = 32'd; 
32'd43829: dataIn1 = 32'd; 
32'd43830: dataIn1 = 32'd; 
32'd43831: dataIn1 = 32'd; 
32'd43832: dataIn1 = 32'd; 
32'd43833: dataIn1 = 32'd; 
32'd43834: dataIn1 = 32'd; 
32'd43835: dataIn1 = 32'd; 
32'd43836: dataIn1 = 32'd; 
32'd43837: dataIn1 = 32'd; 
32'd43838: dataIn1 = 32'd; 
32'd43839: dataIn1 = 32'd; 
32'd43840: dataIn1 = 32'd; 
32'd43841: dataIn1 = 32'd; 
32'd43842: dataIn1 = 32'd; 
32'd43843: dataIn1 = 32'd; 
32'd43844: dataIn1 = 32'd; 
32'd43845: dataIn1 = 32'd; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd37; 
32'd3: dataIn2 = 32'd100; 
32'd4: dataIn2 = 32'd3; 
32'd5: dataIn2 = 32'd58; 
32'd6: dataIn2 = 32'd23; 
32'd7: dataIn2 = 32'd56; 
32'd8: dataIn2 = 32'd30; 
32'd9: dataIn2 = 32'd21; 
32'd10: dataIn2 = 32'd3; 
32'd11: dataIn2 = 32'd7; 
32'd12: dataIn2 = 32'd93; 
32'd13: dataIn2 = 32'd57; 
32'd14: dataIn2 = 32'd57; 
32'd15: dataIn2 = 32'd23; 
32'd16: dataIn2 = 32'd55; 
32'd17: dataIn2 = 32'd96; 
32'd18: dataIn2 = 32'd50; 
32'd19: dataIn2 = 32'd97; 
32'd20: dataIn2 = 32'd86; 
32'd21: dataIn2 = 32'd14; 
32'd22: dataIn2 = 32'd51; 
32'd23: dataIn2 = 32'd49; 
32'd24: dataIn2 = 32'd56; 
32'd25: dataIn2 = 32'd70; 
32'd26: dataIn2 = 32'd96; 
32'd27: dataIn2 = 32'd49; 
32'd28: dataIn2 = 32'd47; 
32'd29: dataIn2 = 32'd61; 
32'd30: dataIn2 = 32'd9; 
32'd31: dataIn2 = 32'd50; 
32'd32: dataIn2 = 32'd46; 
32'd33: dataIn2 = 32'd84; 
32'd34: dataIn2 = 32'd55; 
32'd35: dataIn2 = 32'd66; 
32'd36: dataIn2 = 32'd1; 
32'd37: dataIn2 = 32'd90; 
32'd38: dataIn2 = 32'd9; 
32'd39: dataIn2 = 32'd14; 
32'd40: dataIn2 = 32'd14; 
32'd41: dataIn2 = 32'd43; 
32'd42: dataIn2 = 32'd77; 
32'd43: dataIn2 = 32'd29; 
32'd44: dataIn2 = 32'd54; 
32'd45: dataIn2 = 32'd23; 
32'd46: dataIn2 = 32'd36; 
32'd47: dataIn2 = 32'd8; 
32'd48: dataIn2 = 32'd63; 
32'd49: dataIn2 = 32'd77; 
32'd50: dataIn2 = 32'd15; 
32'd51: dataIn2 = 32'd83; 
32'd52: dataIn2 = 32'd50; 
32'd53: dataIn2 = 32'd22; 
32'd54: dataIn2 = 32'd24; 
32'd55: dataIn2 = 32'd26; 
32'd56: dataIn2 = 32'd65; 
32'd57: dataIn2 = 32'd14; 
32'd58: dataIn2 = 32'd71; 
32'd59: dataIn2 = 32'd75; 
32'd60: dataIn2 = 32'd79; 
32'd61: dataIn2 = 32'd5; 
32'd62: dataIn2 = 32'd100; 
32'd63: dataIn2 = 32'd13; 
32'd64: dataIn2 = 32'd41; 
32'd65: dataIn2 = 32'd6; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd330: dataIn2 = 32'd38; 
32'd331: dataIn2 = 32'd45; 
32'd332: dataIn2 = 32'd52; 
32'd333: dataIn2 = 32'd88; 
32'd334: dataIn2 = 32'd21; 
32'd335: dataIn2 = 32'd56; 
32'd336: dataIn2 = 32'd7; 
32'd337: dataIn2 = 32'd25; 
32'd338: dataIn2 = 32'd67; 
32'd339: dataIn2 = 32'd68; 
32'd340: dataIn2 = 32'd10; 
32'd341: dataIn2 = 32'd31; 
32'd342: dataIn2 = 32'd43; 
32'd343: dataIn2 = 32'd55; 
32'd344: dataIn2 = 32'd45; 
32'd345: dataIn2 = 32'd34; 
32'd346: dataIn2 = 32'd99; 
32'd347: dataIn2 = 32'd58; 
32'd348: dataIn2 = 32'd53; 
32'd349: dataIn2 = 32'd26; 
32'd350: dataIn2 = 32'd52; 
32'd351: dataIn2 = 32'd25; 
32'd352: dataIn2 = 32'd20; 
32'd353: dataIn2 = 32'd95; 
32'd354: dataIn2 = 32'd32; 
32'd355: dataIn2 = 32'd43; 
32'd356: dataIn2 = 32'd83; 
32'd357: dataIn2 = 32'd6; 
32'd358: dataIn2 = 32'd39; 
32'd359: dataIn2 = 32'd62; 
32'd360: dataIn2 = 32'd32; 
32'd361: dataIn2 = 32'd0; 
32'd362: dataIn2 = 32'd54; 
32'd363: dataIn2 = 32'd84; 
32'd364: dataIn2 = 32'd10; 
32'd365: dataIn2 = 32'd96; 
32'd366: dataIn2 = 32'd80; 
32'd367: dataIn2 = 32'd50; 
32'd368: dataIn2 = 32'd47; 
32'd369: dataIn2 = 32'd49; 
32'd370: dataIn2 = 32'd6; 
32'd371: dataIn2 = 32'd33; 
32'd372: dataIn2 = 32'd94; 
32'd373: dataIn2 = 32'd65; 
32'd374: dataIn2 = 32'd81; 
32'd375: dataIn2 = 32'd2; 
32'd376: dataIn2 = 32'd37; 
32'd377: dataIn2 = 32'd77; 
32'd378: dataIn2 = 32'd93; 
32'd379: dataIn2 = 32'd78; 
32'd380: dataIn2 = 32'd42; 
32'd381: dataIn2 = 32'd8; 
32'd382: dataIn2 = 32'd52; 
32'd383: dataIn2 = 32'd47; 
32'd384: dataIn2 = 32'd85; 
32'd385: dataIn2 = 32'd51; 
32'd386: dataIn2 = 32'd1; 
32'd387: dataIn2 = 32'd48; 
32'd388: dataIn2 = 32'd7; 
32'd389: dataIn2 = 32'd94; 
32'd390: dataIn2 = 32'd85; 
32'd391: dataIn2 = 32'd69; 
32'd392: dataIn2 = 32'd59; 
32'd393: dataIn2 = 32'd4; 
32'd394: dataIn2 = 32'd19; 
32'd395: dataIn2 = 32'd7; 
32'd396: dataIn2 = 32'd72; 
32'd397: dataIn2 = 32'd4; 
32'd398: dataIn2 = 32'd65; 
32'd399: dataIn2 = 32'd37; 
32'd400: dataIn2 = 32'd58; 
32'd401: dataIn2 = 32'd90; 
32'd402: dataIn2 = 32'd4; 
32'd403: dataIn2 = 32'd100; 
32'd404: dataIn2 = 32'd84; 
32'd405: dataIn2 = 32'd1; 
32'd406: dataIn2 = 32'd67; 
32'd407: dataIn2 = 32'd61; 
32'd408: dataIn2 = 32'd26; 
32'd409: dataIn2 = 32'd38; 
32'd410: dataIn2 = 32'd47; 
32'd411: dataIn2 = 32'd27; 
32'd412: dataIn2 = 32'd13; 
32'd413: dataIn2 = 32'd92; 
32'd414: dataIn2 = 32'd77; 
32'd415: dataIn2 = 32'd83; 
32'd416: dataIn2 = 32'd46; 
32'd417: dataIn2 = 32'd46; 
32'd418: dataIn2 = 32'd47; 
32'd419: dataIn2 = 32'd39; 
32'd420: dataIn2 = 32'd61; 
32'd421: dataIn2 = 32'd11; 
32'd422: dataIn2 = 32'd40; 
32'd423: dataIn2 = 32'd9; 
32'd424: dataIn2 = 32'd32; 
32'd425: dataIn2 = 32'd65; 
32'd426: dataIn2 = 32'd10; 
32'd427: dataIn2 = 32'd24; 
32'd428: dataIn2 = 32'd9; 
32'd429: dataIn2 = 32'd8; 
32'd430: dataIn2 = 32'd3; 
32'd431: dataIn2 = 32'd89; 
32'd432: dataIn2 = 32'd43; 
32'd433: dataIn2 = 32'd8; 
32'd434: dataIn2 = 32'd68; 
32'd435: dataIn2 = 32'd33; 
32'd436: dataIn2 = 32'd25; 
32'd437: dataIn2 = 32'd86; 
32'd438: dataIn2 = 32'd7; 
32'd439: dataIn2 = 32'd37; 
32'd440: dataIn2 = 32'd78; 
32'd441: dataIn2 = 32'd50; 
32'd442: dataIn2 = 32'd55; 
32'd443: dataIn2 = 32'd63; 
32'd444: dataIn2 = 32'd39; 
32'd445: dataIn2 = 32'd67; 
32'd446: dataIn2 = 32'd18; 
32'd447: dataIn2 = 32'd1; 
32'd448: dataIn2 = 32'd78; 
32'd449: dataIn2 = 32'd85; 
32'd450: dataIn2 = 32'd40; 
32'd451: dataIn2 = 32'd60; 
32'd452: dataIn2 = 32'd49; 
32'd453: dataIn2 = 32'd84; 
32'd454: dataIn2 = 32'd99; 
32'd455: dataIn2 = 32'd92; 
32'd456: dataIn2 = 32'd36; 
32'd457: dataIn2 = 32'd20; 
32'd458: dataIn2 = 32'd95; 
32'd459: dataIn2 = 32'd17; 
32'd460: dataIn2 = 32'd49; 
32'd461: dataIn2 = 32'd97; 
32'd462: dataIn2 = 32'd76; 
32'd463: dataIn2 = 32'd79; 
32'd464: dataIn2 = 32'd16; 
32'd465: dataIn2 = 32'd60; 
32'd466: dataIn2 = 32'd82; 
32'd467: dataIn2 = 32'd85; 
32'd468: dataIn2 = 32'd55; 
32'd469: dataIn2 = 32'd72; 
32'd470: dataIn2 = 32'd96; 
32'd471: dataIn2 = 32'd80; 
32'd472: dataIn2 = 32'd72; 
32'd473: dataIn2 = 32'd59; 
32'd474: dataIn2 = 32'd18; 
32'd475: dataIn2 = 32'd60; 
32'd476: dataIn2 = 32'd52; 
32'd477: dataIn2 = 32'd87; 
32'd478: dataIn2 = 32'd74; 
32'd479: dataIn2 = 32'd98; 
32'd480: dataIn2 = 32'd17; 
32'd481: dataIn2 = 32'd60; 
32'd482: dataIn2 = 32'd71; 
32'd483: dataIn2 = 32'd80; 
32'd484: dataIn2 = 32'd59; 
32'd485: dataIn2 = 32'd55; 
32'd486: dataIn2 = 32'd9; 
32'd487: dataIn2 = 32'd59; 
32'd488: dataIn2 = 32'd14; 
32'd489: dataIn2 = 32'd22; 
32'd490: dataIn2 = 32'd71; 
32'd491: dataIn2 = 32'd93; 
32'd492: dataIn2 = 32'd58; 
32'd493: dataIn2 = 32'd55; 
32'd494: dataIn2 = 32'd62; 
32'd495: dataIn2 = 32'd6; 
32'd496: dataIn2 = 32'd71; 
32'd497: dataIn2 = 32'd29; 
32'd498: dataIn2 = 32'd39; 
32'd499: dataIn2 = 32'd22; 
32'd500: dataIn2 = 32'd48; 
32'd501: dataIn2 = 32'd20; 
32'd502: dataIn2 = 32'd7; 
32'd503: dataIn2 = 32'd58; 
32'd504: dataIn2 = 32'd87; 
32'd505: dataIn2 = 32'd30; 
32'd506: dataIn2 = 32'd66; 
32'd507: dataIn2 = 32'd47; 
32'd508: dataIn2 = 32'd49; 
32'd509: dataIn2 = 32'd86; 
32'd510: dataIn2 = 32'd43; 
32'd511: dataIn2 = 32'd78; 
32'd512: dataIn2 = 32'd50; 
32'd513: dataIn2 = 32'd59; 
32'd514: dataIn2 = 32'd36; 
32'd515: dataIn2 = 32'd5; 
32'd516: dataIn2 = 32'd17; 
32'd517: dataIn2 = 32'd53; 
32'd518: dataIn2 = 32'd33; 
32'd519: dataIn2 = 32'd100; 
32'd520: dataIn2 = 32'd70; 
32'd521: dataIn2 = 32'd48; 
32'd522: dataIn2 = 32'd76; 
32'd523: dataIn2 = 32'd72; 
32'd524: dataIn2 = 32'd60; 
32'd525: dataIn2 = 32'd87; 
32'd526: dataIn2 = 32'd28; 
32'd527: dataIn2 = 32'd48; 
32'd528: dataIn2 = 32'd55; 
32'd529: dataIn2 = 32'd57; 
32'd530: dataIn2 = 32'd60; 
32'd531: dataIn2 = 32'd61; 
32'd532: dataIn2 = 32'd38; 
32'd533: dataIn2 = 32'd9; 
32'd534: dataIn2 = 32'd50; 
32'd535: dataIn2 = 32'd64; 
32'd536: dataIn2 = 32'd92; 
32'd537: dataIn2 = 32'd84; 
32'd538: dataIn2 = 32'd65; 
32'd539: dataIn2 = 32'd97; 
32'd540: dataIn2 = 32'd74; 
32'd541: dataIn2 = 32'd71; 
32'd542: dataIn2 = 32'd5; 
32'd543: dataIn2 = 32'd78; 
32'd544: dataIn2 = 32'd79; 
32'd545: dataIn2 = 32'd47; 
32'd546: dataIn2 = 32'd39; 
32'd547: dataIn2 = 32'd80; 
32'd548: dataIn2 = 32'd53; 
32'd549: dataIn2 = 32'd65; 
32'd550: dataIn2 = 32'd72; 
32'd551: dataIn2 = 32'd74; 
32'd552: dataIn2 = 32'd80; 
32'd553: dataIn2 = 32'd10; 
32'd554: dataIn2 = 32'd43; 
32'd555: dataIn2 = 32'd84; 
32'd556: dataIn2 = 32'd19; 
32'd557: dataIn2 = 32'd28; 
32'd558: dataIn2 = 32'd44; 
32'd559: dataIn2 = 32'd47; 
32'd560: dataIn2 = 32'd91; 
32'd561: dataIn2 = 32'd38; 
32'd562: dataIn2 = 32'd47; 
32'd563: dataIn2 = 32'd69; 
32'd564: dataIn2 = 32'd66; 
32'd565: dataIn2 = 32'd71; 
32'd566: dataIn2 = 32'd60; 
32'd567: dataIn2 = 32'd52; 
32'd568: dataIn2 = 32'd46; 
32'd569: dataIn2 = 32'd85; 
32'd570: dataIn2 = 32'd39; 
32'd571: dataIn2 = 32'd95; 
32'd572: dataIn2 = 32'd95; 
32'd573: dataIn2 = 32'd44; 
32'd574: dataIn2 = 32'd6; 
32'd575: dataIn2 = 32'd27; 
32'd576: dataIn2 = 32'd37; 
32'd577: dataIn2 = 32'd86; 
32'd578: dataIn2 = 32'd55; 
32'd579: dataIn2 = 32'd91; 
32'd580: dataIn2 = 32'd87; 
32'd581: dataIn2 = 32'd2; 
32'd582: dataIn2 = 32'd78; 
32'd583: dataIn2 = 32'd19; 
32'd584: dataIn2 = 32'd88; 
32'd585: dataIn2 = 32'd80; 
32'd586: dataIn2 = 32'd98; 
32'd587: dataIn2 = 32'd95; 
32'd588: dataIn2 = 32'd29; 
32'd589: dataIn2 = 32'd19; 
32'd590: dataIn2 = 32'd73; 
32'd591: dataIn2 = 32'd76; 
32'd592: dataIn2 = 32'd89; 
32'd593: dataIn2 = 32'd73; 
32'd594: dataIn2 = 32'd25; 
32'd595: dataIn2 = 32'd27; 
32'd596: dataIn2 = 32'd67; 
32'd597: dataIn2 = 32'd56; 
32'd598: dataIn2 = 32'd54; 
32'd599: dataIn2 = 32'd40; 
32'd600: dataIn2 = 32'd60; 
32'd601: dataIn2 = 32'd59; 
32'd602: dataIn2 = 32'd43; 
32'd603: dataIn2 = 32'd93; 
32'd604: dataIn2 = 32'd73; 
32'd605: dataIn2 = 32'd54; 
32'd606: dataIn2 = 32'd14; 
32'd607: dataIn2 = 32'd1; 
32'd608: dataIn2 = 32'd15; 
32'd609: dataIn2 = 32'd95; 
32'd610: dataIn2 = 32'd98; 
32'd611: dataIn2 = 32'd22; 
32'd612: dataIn2 = 32'd29; 
32'd613: dataIn2 = 32'd96; 
32'd614: dataIn2 = 32'd52; 
32'd615: dataIn2 = 32'd71; 
32'd616: dataIn2 = 32'd78; 
32'd617: dataIn2 = 32'd78; 
32'd618: dataIn2 = 32'd25; 
32'd619: dataIn2 = 32'd31; 
32'd620: dataIn2 = 32'd2; 
32'd621: dataIn2 = 32'd43; 
32'd622: dataIn2 = 32'd46; 
32'd623: dataIn2 = 32'd23; 
32'd624: dataIn2 = 32'd26; 
32'd625: dataIn2 = 32'd8; 
32'd626: dataIn2 = 32'd88; 
32'd627: dataIn2 = 32'd38; 
32'd628: dataIn2 = 32'd15; 
32'd629: dataIn2 = 32'd88; 
32'd630: dataIn2 = 32'd25; 
32'd631: dataIn2 = 32'd20; 
32'd632: dataIn2 = 32'd49; 
32'd633: dataIn2 = 32'd36; 
32'd634: dataIn2 = 32'd84; 
32'd635: dataIn2 = 32'd32; 
32'd636: dataIn2 = 32'd0; 
32'd637: dataIn2 = 32'd79; 
32'd638: dataIn2 = 32'd23; 
32'd639: dataIn2 = 32'd92; 
32'd640: dataIn2 = 32'd10; 
32'd641: dataIn2 = 32'd5; 
32'd642: dataIn2 = 32'd35; 
32'd643: dataIn2 = 32'd23; 
32'd644: dataIn2 = 32'd56; 
32'd645: dataIn2 = 32'd18; 
32'd646: dataIn2 = 32'd80; 
32'd647: dataIn2 = 32'd18; 
32'd648: dataIn2 = 32'd90; 
32'd649: dataIn2 = 32'd6; 
32'd650: dataIn2 = 32'd31; 
32'd651: dataIn2 = 32'd4; 
32'd652: dataIn2 = 32'd32; 
32'd653: dataIn2 = 32'd19; 
32'd654: dataIn2 = 32'd0; 
32'd655: dataIn2 = 32'd84; 
32'd656: dataIn2 = 32'd37; 
32'd657: dataIn2 = 32'd54; 
32'd658: dataIn2 = 32'd43; 
32'd659: dataIn2 = 32'd17; 
32'd660: dataIn2 = 32'd25; 
32'd661: dataIn2 = 32'd7; 
32'd662: dataIn2 = 32'd15; 
32'd663: dataIn2 = 32'd94; 
32'd664: dataIn2 = 32'd7; 
32'd665: dataIn2 = 32'd60; 
32'd666: dataIn2 = 32'd17; 
32'd667: dataIn2 = 32'd1; 
32'd668: dataIn2 = 32'd9; 
32'd669: dataIn2 = 32'd24; 
32'd670: dataIn2 = 32'd96; 
32'd671: dataIn2 = 32'd57; 
32'd672: dataIn2 = 32'd83; 
32'd673: dataIn2 = 32'd85; 
32'd674: dataIn2 = 32'd5; 
32'd675: dataIn2 = 32'd47; 
32'd676: dataIn2 = 32'd76; 
32'd677: dataIn2 = 32'd36; 
32'd678: dataIn2 = 32'd10; 
32'd679: dataIn2 = 32'd93; 
32'd680: dataIn2 = 32'd8; 
32'd681: dataIn2 = 32'd0; 
32'd682: dataIn2 = 32'd47; 
32'd683: dataIn2 = 32'd53; 
32'd684: dataIn2 = 32'd69; 
32'd685: dataIn2 = 32'd12; 
32'd686: dataIn2 = 32'd57; 
32'd687: dataIn2 = 32'd7; 
32'd688: dataIn2 = 32'd73; 
32'd689: dataIn2 = 32'd85; 
32'd690: dataIn2 = 32'd4; 
32'd691: dataIn2 = 32'd45; 
32'd692: dataIn2 = 32'd40; 
32'd693: dataIn2 = 32'd15; 
32'd694: dataIn2 = 32'd11; 
32'd695: dataIn2 = 32'd97; 
32'd696: dataIn2 = 32'd88; 
32'd697: dataIn2 = 32'd69; 
32'd698: dataIn2 = 32'd97; 
32'd699: dataIn2 = 32'd25; 
32'd700: dataIn2 = 32'd16; 
32'd701: dataIn2 = 32'd5; 
32'd702: dataIn2 = 32'd51; 
32'd703: dataIn2 = 32'd26; 
32'd704: dataIn2 = 32'd4; 
32'd705: dataIn2 = 32'd54; 
32'd706: dataIn2 = 32'd54; 
32'd707: dataIn2 = 32'd90; 
32'd708: dataIn2 = 32'd57; 
32'd709: dataIn2 = 32'd47; 
32'd710: dataIn2 = 32'd24; 
32'd711: dataIn2 = 32'd70; 
32'd712: dataIn2 = 32'd81; 
32'd713: dataIn2 = 32'd39; 
32'd714: dataIn2 = 32'd82; 
32'd715: dataIn2 = 32'd4; 
32'd716: dataIn2 = 32'd47; 
32'd717: dataIn2 = 32'd31; 
32'd718: dataIn2 = 32'd67; 
32'd719: dataIn2 = 32'd81; 
32'd720: dataIn2 = 32'd51; 
32'd721: dataIn2 = 32'd80; 
32'd722: dataIn2 = 32'd29; 
32'd723: dataIn2 = 32'd39; 
32'd724: dataIn2 = 32'd20; 
32'd725: dataIn2 = 32'd82; 
32'd726: dataIn2 = 32'd73; 
32'd727: dataIn2 = 32'd88; 
32'd728: dataIn2 = 32'd1; 
32'd729: dataIn2 = 32'd69; 
32'd730: dataIn2 = 32'd25; 
32'd731: dataIn2 = 32'd5; 
32'd732: dataIn2 = 32'd44; 
32'd733: dataIn2 = 32'd42; 
32'd734: dataIn2 = 32'd100; 
32'd735: dataIn2 = 32'd40; 
32'd736: dataIn2 = 32'd20; 
32'd737: dataIn2 = 32'd9; 
32'd738: dataIn2 = 32'd71; 
32'd739: dataIn2 = 32'd75; 
32'd740: dataIn2 = 32'd77; 
32'd741: dataIn2 = 32'd20; 
32'd742: dataIn2 = 32'd60; 
32'd743: dataIn2 = 32'd35; 
32'd744: dataIn2 = 32'd1; 
32'd745: dataIn2 = 32'd29; 
32'd746: dataIn2 = 32'd67; 
32'd747: dataIn2 = 32'd35; 
32'd748: dataIn2 = 32'd8; 
32'd749: dataIn2 = 32'd80; 
32'd750: dataIn2 = 32'd53; 
32'd751: dataIn2 = 32'd84; 
32'd752: dataIn2 = 32'd29; 
32'd753: dataIn2 = 32'd46; 
32'd754: dataIn2 = 32'd86; 
32'd755: dataIn2 = 32'd58; 
32'd756: dataIn2 = 32'd22; 
32'd757: dataIn2 = 32'd43; 
32'd758: dataIn2 = 32'd17; 
32'd759: dataIn2 = 32'd44; 
32'd760: dataIn2 = 32'd79; 
32'd761: dataIn2 = 32'd50; 
32'd762: dataIn2 = 32'd21; 
32'd763: dataIn2 = 32'd50; 
32'd764: dataIn2 = 32'd98; 
32'd765: dataIn2 = 32'd69; 
32'd766: dataIn2 = 32'd98; 
32'd767: dataIn2 = 32'd82; 
32'd768: dataIn2 = 32'd37; 
32'd769: dataIn2 = 32'd4; 
32'd770: dataIn2 = 32'd76; 
32'd771: dataIn2 = 32'd87; 
32'd772: dataIn2 = 32'd40; 
32'd773: dataIn2 = 32'd1; 
32'd774: dataIn2 = 32'd68; 
32'd775: dataIn2 = 32'd57; 
32'd776: dataIn2 = 32'd6; 
32'd777: dataIn2 = 32'd29; 
32'd778: dataIn2 = 32'd39; 
32'd779: dataIn2 = 32'd45; 
32'd780: dataIn2 = 32'd18; 
32'd781: dataIn2 = 32'd55; 
32'd782: dataIn2 = 32'd96; 
32'd783: dataIn2 = 32'd48; 
32'd784: dataIn2 = 32'd17; 
32'd785: dataIn2 = 32'd65; 
32'd786: dataIn2 = 32'd35; 
32'd787: dataIn2 = 32'd79; 
32'd788: dataIn2 = 32'd53; 
32'd789: dataIn2 = 32'd67; 
32'd790: dataIn2 = 32'd75; 
32'd791: dataIn2 = 32'd48; 
32'd792: dataIn2 = 32'd66; 
32'd793: dataIn2 = 32'd92; 
32'd794: dataIn2 = 32'd75; 
32'd795: dataIn2 = 32'd21; 
32'd796: dataIn2 = 32'd81; 
32'd797: dataIn2 = 32'd26; 
32'd798: dataIn2 = 32'd36; 
32'd799: dataIn2 = 32'd53; 
32'd800: dataIn2 = 32'd78; 
32'd801: dataIn2 = 32'd100; 
32'd802: dataIn2 = 32'd0; 
32'd803: dataIn2 = 32'd0; 
32'd804: dataIn2 = 32'd73; 
32'd805: dataIn2 = 32'd54; 
32'd806: dataIn2 = 32'd77; 
32'd807: dataIn2 = 32'd91; 
32'd808: dataIn2 = 32'd5; 
32'd809: dataIn2 = 32'd21; 
32'd810: dataIn2 = 32'd28; 
32'd811: dataIn2 = 32'd9; 
32'd812: dataIn2 = 32'd71; 
32'd813: dataIn2 = 32'd53; 
32'd814: dataIn2 = 32'd71; 
32'd815: dataIn2 = 32'd42; 
32'd816: dataIn2 = 32'd99; 
32'd817: dataIn2 = 32'd21; 
32'd818: dataIn2 = 32'd43; 
32'd819: dataIn2 = 32'd54; 
32'd820: dataIn2 = 32'd44; 
32'd821: dataIn2 = 32'd29; 
32'd822: dataIn2 = 32'd54; 
32'd823: dataIn2 = 32'd79; 
32'd824: dataIn2 = 32'd55; 
32'd825: dataIn2 = 32'd17; 
32'd826: dataIn2 = 32'd34; 
32'd827: dataIn2 = 32'd27; 
32'd828: dataIn2 = 32'd9; 
32'd829: dataIn2 = 32'd34; 
32'd830: dataIn2 = 32'd97; 
32'd831: dataIn2 = 32'd73; 
32'd832: dataIn2 = 32'd59; 
32'd833: dataIn2 = 32'd48; 
32'd834: dataIn2 = 32'd47; 
32'd835: dataIn2 = 32'd52; 
32'd836: dataIn2 = 32'd12; 
32'd837: dataIn2 = 32'd91; 
32'd838: dataIn2 = 32'd23; 
32'd839: dataIn2 = 32'd100; 
32'd840: dataIn2 = 32'd68; 
32'd841: dataIn2 = 32'd62; 
32'd842: dataIn2 = 32'd5; 
32'd843: dataIn2 = 32'd90; 
32'd844: dataIn2 = 32'd47; 
32'd845: dataIn2 = 32'd78; 
32'd846: dataIn2 = 32'd16; 
32'd847: dataIn2 = 32'd91; 
32'd848: dataIn2 = 32'd21; 
32'd849: dataIn2 = 32'd25; 
32'd850: dataIn2 = 32'd62; 
32'd851: dataIn2 = 32'd5; 
32'd852: dataIn2 = 32'd93; 
32'd853: dataIn2 = 32'd31; 
32'd854: dataIn2 = 32'd61; 
32'd855: dataIn2 = 32'd13; 
32'd856: dataIn2 = 32'd75; 
32'd857: dataIn2 = 32'd90; 
32'd858: dataIn2 = 32'd90; 
32'd859: dataIn2 = 32'd56; 
32'd860: dataIn2 = 32'd55; 
32'd861: dataIn2 = 32'd61; 
32'd862: dataIn2 = 32'd33; 
32'd863: dataIn2 = 32'd11; 
32'd864: dataIn2 = 32'd11; 
32'd865: dataIn2 = 32'd11; 
32'd866: dataIn2 = 32'd9; 
32'd867: dataIn2 = 32'd38; 
32'd868: dataIn2 = 32'd48; 
32'd869: dataIn2 = 32'd49; 
32'd870: dataIn2 = 32'd10; 
32'd871: dataIn2 = 32'd1; 
32'd872: dataIn2 = 32'd2; 
32'd873: dataIn2 = 32'd79; 
32'd874: dataIn2 = 32'd27; 
32'd875: dataIn2 = 32'd85; 
32'd876: dataIn2 = 32'd26; 
32'd877: dataIn2 = 32'd10; 
32'd878: dataIn2 = 32'd4; 
32'd879: dataIn2 = 32'd73; 
32'd880: dataIn2 = 32'd83; 
32'd881: dataIn2 = 32'd86; 
32'd882: dataIn2 = 32'd3; 
32'd883: dataIn2 = 32'd0; 
32'd884: dataIn2 = 32'd1; 
32'd885: dataIn2 = 32'd35; 
32'd886: dataIn2 = 32'd67; 
32'd887: dataIn2 = 32'd26; 
32'd888: dataIn2 = 32'd53; 
32'd889: dataIn2 = 32'd30; 
32'd890: dataIn2 = 32'd77; 
32'd891: dataIn2 = 32'd1; 
32'd892: dataIn2 = 32'd16; 
32'd893: dataIn2 = 32'd35; 
32'd894: dataIn2 = 32'd31; 
32'd895: dataIn2 = 32'd45; 
32'd896: dataIn2 = 32'd93; 
32'd897: dataIn2 = 32'd15; 
32'd898: dataIn2 = 32'd63; 
32'd899: dataIn2 = 32'd46; 
32'd900: dataIn2 = 32'd8; 
32'd901: dataIn2 = 32'd55; 
32'd902: dataIn2 = 32'd63; 
32'd903: dataIn2 = 32'd17; 
32'd904: dataIn2 = 32'd80; 
32'd905: dataIn2 = 32'd44; 
32'd906: dataIn2 = 32'd2; 
32'd907: dataIn2 = 32'd44; 
32'd908: dataIn2 = 32'd67; 
32'd909: dataIn2 = 32'd20; 
32'd910: dataIn2 = 32'd22; 
32'd911: dataIn2 = 32'd70; 
32'd912: dataIn2 = 32'd18; 
32'd913: dataIn2 = 32'd92; 
32'd914: dataIn2 = 32'd85; 
32'd915: dataIn2 = 32'd31; 
32'd916: dataIn2 = 32'd43; 
32'd917: dataIn2 = 32'd33; 
32'd918: dataIn2 = 32'd94; 
32'd919: dataIn2 = 32'd79; 
32'd920: dataIn2 = 32'd41; 
32'd921: dataIn2 = 32'd95; 
32'd922: dataIn2 = 32'd79; 
32'd923: dataIn2 = 32'd83; 
32'd924: dataIn2 = 32'd97; 
32'd925: dataIn2 = 32'd62; 
32'd926: dataIn2 = 32'd95; 
32'd927: dataIn2 = 32'd21; 
32'd928: dataIn2 = 32'd13; 
32'd929: dataIn2 = 32'd81; 
32'd930: dataIn2 = 32'd24; 
32'd931: dataIn2 = 32'd15; 
32'd932: dataIn2 = 32'd60; 
32'd933: dataIn2 = 32'd91; 
32'd934: dataIn2 = 32'd60; 
32'd935: dataIn2 = 32'd38; 
32'd936: dataIn2 = 32'd45; 
32'd937: dataIn2 = 32'd43; 
32'd938: dataIn2 = 32'd59; 
32'd939: dataIn2 = 32'd24; 
32'd940: dataIn2 = 32'd40; 
32'd941: dataIn2 = 32'd87; 
32'd942: dataIn2 = 32'd73; 
32'd943: dataIn2 = 32'd43; 
32'd944: dataIn2 = 32'd33; 
32'd945: dataIn2 = 32'd71; 
32'd946: dataIn2 = 32'd12; 
32'd947: dataIn2 = 32'd84; 
32'd948: dataIn2 = 32'd53; 
32'd949: dataIn2 = 32'd2; 
32'd950: dataIn2 = 32'd91; 
32'd951: dataIn2 = 32'd23; 
32'd952: dataIn2 = 32'd55; 
32'd953: dataIn2 = 32'd51; 
32'd954: dataIn2 = 32'd74; 
32'd955: dataIn2 = 32'd48; 
32'd956: dataIn2 = 32'd15; 
32'd957: dataIn2 = 32'd73; 
32'd958: dataIn2 = 32'd54; 
32'd959: dataIn2 = 32'd48; 
32'd960: dataIn2 = 32'd98; 
32'd961: dataIn2 = 32'd53; 
32'd962: dataIn2 = 32'd7; 
32'd963: dataIn2 = 32'd57; 
32'd964: dataIn2 = 32'd45; 
32'd965: dataIn2 = 32'd91; 
32'd966: dataIn2 = 32'd25; 
32'd967: dataIn2 = 32'd80; 
32'd968: dataIn2 = 32'd89; 
32'd969: dataIn2 = 32'd31; 
32'd970: dataIn2 = 32'd99; 
32'd971: dataIn2 = 32'd86; 
32'd972: dataIn2 = 32'd28; 
32'd973: dataIn2 = 32'd35; 
32'd974: dataIn2 = 32'd31; 
32'd975: dataIn2 = 32'd7; 
32'd976: dataIn2 = 32'd6; 
32'd977: dataIn2 = 32'd79; 
32'd978: dataIn2 = 32'd57; 
32'd979: dataIn2 = 32'd62; 
32'd980: dataIn2 = 32'd93; 
32'd981: dataIn2 = 32'd18; 
32'd982: dataIn2 = 32'd9; 
32'd983: dataIn2 = 32'd65; 
32'd984: dataIn2 = 32'd37; 
32'd985: dataIn2 = 32'd7; 
32'd986: dataIn2 = 32'd49; 
32'd987: dataIn2 = 32'd35; 
32'd988: dataIn2 = 32'd42; 
32'd989: dataIn2 = 32'd100; 
32'd990: dataIn2 = 32'd36; 
32'd991: dataIn2 = 32'd96; 
32'd992: dataIn2 = 32'd1; 
32'd993: dataIn2 = 32'd22; 
32'd994: dataIn2 = 32'd68; 
32'd995: dataIn2 = 32'd73; 
32'd996: dataIn2 = 32'd83; 
32'd997: dataIn2 = 32'd22; 
32'd998: dataIn2 = 32'd98; 
32'd999: dataIn2 = 32'd41; 
32'd1000: dataIn2 = 32'd76; 
32'd1001: dataIn2 = 32'd30; 
32'd1002: dataIn2 = 32'd62; 
32'd1003: dataIn2 = 32'd63; 
32'd1004: dataIn2 = 32'd95; 
32'd1005: dataIn2 = 32'd71; 
32'd1006: dataIn2 = 32'd58; 
32'd1007: dataIn2 = 32'd19; 
32'd1008: dataIn2 = 32'd66; 
32'd1009: dataIn2 = 32'd55; 
32'd1010: dataIn2 = 32'd33; 
32'd1011: dataIn2 = 32'd67; 
32'd1012: dataIn2 = 32'd51; 
32'd1013: dataIn2 = 32'd64; 
32'd1014: dataIn2 = 32'd11; 
32'd1015: dataIn2 = 32'd42; 
32'd1016: dataIn2 = 32'd13; 
32'd1017: dataIn2 = 32'd38; 
32'd1018: dataIn2 = 32'd53; 
32'd1019: dataIn2 = 32'd35; 
32'd1020: dataIn2 = 32'd68; 
32'd1021: dataIn2 = 32'd50; 
32'd1022: dataIn2 = 32'd30; 
32'd1023: dataIn2 = 32'd22; 
32'd1024: dataIn2 = 32'd74; 
32'd1025: dataIn2 = 32'd41; 
32'd1026: dataIn2 = 32'd96; 
32'd1027: dataIn2 = 32'd22; 
32'd1028: dataIn2 = 32'd86; 
32'd1029: dataIn2 = 32'd7; 
32'd1030: dataIn2 = 32'd63; 
32'd1031: dataIn2 = 32'd81; 
32'd1032: dataIn2 = 32'd11; 
32'd1033: dataIn2 = 32'd93; 
32'd1034: dataIn2 = 32'd90; 
32'd1035: dataIn2 = 32'd77; 
32'd1036: dataIn2 = 32'd97; 
32'd1037: dataIn2 = 32'd95; 
32'd1038: dataIn2 = 32'd46; 
32'd1039: dataIn2 = 32'd22; 
32'd1040: dataIn2 = 32'd72; 
32'd1041: dataIn2 = 32'd95; 
32'd1042: dataIn2 = 32'd18; 
32'd1043: dataIn2 = 32'd4; 
32'd1044: dataIn2 = 32'd19; 
32'd1045: dataIn2 = 32'd90; 
32'd1046: dataIn2 = 32'd94; 
32'd1047: dataIn2 = 32'd12; 
32'd1048: dataIn2 = 32'd20; 
32'd1049: dataIn2 = 32'd87; 
32'd1050: dataIn2 = 32'd8; 
32'd1051: dataIn2 = 32'd10; 
32'd1052: dataIn2 = 32'd5; 
32'd1053: dataIn2 = 32'd66; 
32'd1054: dataIn2 = 32'd94; 
32'd1055: dataIn2 = 32'd80; 
32'd1056: dataIn2 = 32'd72; 
32'd1057: dataIn2 = 32'd53; 
32'd1058: dataIn2 = 32'd20; 
32'd1059: dataIn2 = 32'd30; 
32'd1060: dataIn2 = 32'd51; 
32'd1061: dataIn2 = 32'd31; 
32'd1062: dataIn2 = 32'd10; 
32'd1063: dataIn2 = 32'd24; 
32'd1064: dataIn2 = 32'd12; 
32'd1065: dataIn2 = 32'd46; 
32'd1066: dataIn2 = 32'd8; 
32'd1067: dataIn2 = 32'd73; 
32'd1068: dataIn2 = 32'd35; 
32'd1069: dataIn2 = 32'd11; 
32'd1070: dataIn2 = 32'd20; 
32'd1071: dataIn2 = 32'd68; 
32'd1072: dataIn2 = 32'd24; 
32'd1073: dataIn2 = 32'd67; 
32'd1074: dataIn2 = 32'd8; 
32'd1075: dataIn2 = 32'd85; 
32'd1076: dataIn2 = 32'd67; 
32'd1077: dataIn2 = 32'd43; 
32'd1078: dataIn2 = 32'd31; 
32'd1079: dataIn2 = 32'd51; 
32'd1080: dataIn2 = 32'd90; 
32'd1081: dataIn2 = 32'd85; 
32'd1082: dataIn2 = 32'd46; 
32'd1083: dataIn2 = 32'd25; 
32'd1084: dataIn2 = 32'd99; 
32'd1085: dataIn2 = 32'd21; 
32'd1086: dataIn2 = 32'd77; 
32'd1087: dataIn2 = 32'd70; 
32'd1088: dataIn2 = 32'd27; 
32'd1089: dataIn2 = 32'd93; 
32'd1090: dataIn2 = 32'd52; 
32'd1091: dataIn2 = 32'd69; 
32'd1092: dataIn2 = 32'd68; 
32'd1093: dataIn2 = 32'd33; 
32'd1094: dataIn2 = 32'd13; 
32'd1095: dataIn2 = 32'd25; 
32'd1096: dataIn2 = 32'd49; 
32'd1097: dataIn2 = 32'd43; 
32'd1098: dataIn2 = 32'd9; 
32'd1099: dataIn2 = 32'd27; 
32'd1100: dataIn2 = 32'd78; 
32'd1101: dataIn2 = 32'd23; 
32'd1102: dataIn2 = 32'd75; 
32'd1103: dataIn2 = 32'd68; 
32'd1104: dataIn2 = 32'd95; 
32'd1105: dataIn2 = 32'd13; 
32'd1106: dataIn2 = 32'd83; 
32'd1107: dataIn2 = 32'd62; 
32'd1108: dataIn2 = 32'd90; 
32'd1109: dataIn2 = 32'd3; 
32'd1110: dataIn2 = 32'd49; 
32'd1111: dataIn2 = 32'd71; 
32'd1112: dataIn2 = 32'd5; 
32'd1113: dataIn2 = 32'd15; 
32'd1114: dataIn2 = 32'd43; 
32'd1115: dataIn2 = 32'd68; 
32'd1116: dataIn2 = 32'd10; 
32'd1117: dataIn2 = 32'd80; 
32'd1118: dataIn2 = 32'd0; 
32'd1119: dataIn2 = 32'd91; 
32'd1120: dataIn2 = 32'd99; 
32'd1121: dataIn2 = 32'd58; 
32'd1122: dataIn2 = 32'd49; 
32'd1123: dataIn2 = 32'd42; 
32'd1124: dataIn2 = 32'd47; 
32'd1125: dataIn2 = 32'd32; 
32'd1126: dataIn2 = 32'd70; 
32'd1127: dataIn2 = 32'd32; 
32'd1128: dataIn2 = 32'd76; 
32'd1129: dataIn2 = 32'd79; 
32'd1130: dataIn2 = 32'd11; 
32'd1131: dataIn2 = 32'd82; 
32'd1132: dataIn2 = 32'd39; 
32'd1133: dataIn2 = 32'd45; 
32'd1134: dataIn2 = 32'd79; 
32'd1135: dataIn2 = 32'd15; 
32'd1136: dataIn2 = 32'd94; 
32'd1137: dataIn2 = 32'd20; 
32'd1138: dataIn2 = 32'd41; 
32'd1139: dataIn2 = 32'd41; 
32'd1140: dataIn2 = 32'd13; 
32'd1141: dataIn2 = 32'd54; 
32'd1142: dataIn2 = 32'd83; 
32'd1143: dataIn2 = 32'd60; 
32'd1144: dataIn2 = 32'd31; 
32'd1145: dataIn2 = 32'd61; 
32'd1146: dataIn2 = 32'd90; 
32'd1147: dataIn2 = 32'd13; 
32'd1148: dataIn2 = 32'd69; 
32'd1149: dataIn2 = 32'd39; 
32'd1150: dataIn2 = 32'd76; 
32'd1151: dataIn2 = 32'd46; 
32'd1152: dataIn2 = 32'd33; 
32'd1153: dataIn2 = 32'd36; 
32'd1154: dataIn2 = 32'd96; 
32'd1155: dataIn2 = 32'd13; 
32'd1156: dataIn2 = 32'd74; 
32'd1157: dataIn2 = 32'd56; 
32'd1158: dataIn2 = 32'd89; 
32'd1159: dataIn2 = 32'd15; 
32'd1160: dataIn2 = 32'd44; 
32'd1161: dataIn2 = 32'd99; 
32'd1162: dataIn2 = 32'd21; 
32'd1163: dataIn2 = 32'd2; 
32'd1164: dataIn2 = 32'd88; 
32'd1165: dataIn2 = 32'd83; 
32'd1166: dataIn2 = 32'd34; 
32'd1167: dataIn2 = 32'd61; 
32'd1168: dataIn2 = 32'd22; 
32'd1169: dataIn2 = 32'd71; 
32'd1170: dataIn2 = 32'd99; 
32'd1171: dataIn2 = 32'd89; 
32'd1172: dataIn2 = 32'd33; 
32'd1173: dataIn2 = 32'd50; 
32'd1174: dataIn2 = 32'd42; 
32'd1175: dataIn2 = 32'd16; 
32'd1176: dataIn2 = 32'd84; 
32'd1177: dataIn2 = 32'd33; 
32'd1178: dataIn2 = 32'd46; 
32'd1179: dataIn2 = 32'd71; 
32'd1180: dataIn2 = 32'd81; 
32'd1181: dataIn2 = 32'd83; 
32'd1182: dataIn2 = 32'd48; 
32'd1183: dataIn2 = 32'd20; 
32'd1184: dataIn2 = 32'd41; 
32'd1185: dataIn2 = 32'd11; 
32'd1186: dataIn2 = 32'd82; 
32'd1187: dataIn2 = 32'd15; 
32'd1188: dataIn2 = 32'd94; 
32'd1189: dataIn2 = 32'd85; 
32'd1190: dataIn2 = 32'd50; 
32'd1191: dataIn2 = 32'd30; 
32'd1192: dataIn2 = 32'd81; 
32'd1193: dataIn2 = 32'd6; 
32'd1194: dataIn2 = 32'd41; 
32'd1195: dataIn2 = 32'd70; 
32'd1196: dataIn2 = 32'd65; 
32'd1197: dataIn2 = 32'd46; 
32'd1198: dataIn2 = 32'd44; 
32'd1199: dataIn2 = 32'd87; 
32'd1200: dataIn2 = 32'd84; 
32'd1201: dataIn2 = 32'd75; 
32'd1202: dataIn2 = 32'd28; 
32'd1203: dataIn2 = 32'd25; 
32'd1204: dataIn2 = 32'd27; 
32'd1205: dataIn2 = 32'd70; 
32'd1206: dataIn2 = 32'd80; 
32'd1207: dataIn2 = 32'd79; 
32'd1208: dataIn2 = 32'd100; 
32'd1209: dataIn2 = 32'd6; 
32'd1210: dataIn2 = 32'd14; 
32'd1211: dataIn2 = 32'd48; 
32'd1212: dataIn2 = 32'd95; 
32'd1213: dataIn2 = 32'd95; 
32'd1214: dataIn2 = 32'd11; 
32'd1215: dataIn2 = 32'd98; 
32'd1216: dataIn2 = 32'd75; 
32'd1217: dataIn2 = 32'd15; 
32'd1218: dataIn2 = 32'd50; 
32'd1219: dataIn2 = 32'd7; 
32'd1220: dataIn2 = 32'd5; 
32'd1221: dataIn2 = 32'd75; 
32'd1222: dataIn2 = 32'd90; 
32'd1223: dataIn2 = 32'd30; 
32'd1224: dataIn2 = 32'd18; 
32'd1225: dataIn2 = 32'd47; 
32'd1226: dataIn2 = 32'd19; 
32'd1227: dataIn2 = 32'd37; 
32'd1228: dataIn2 = 32'd36; 
32'd1229: dataIn2 = 32'd2; 
32'd1230: dataIn2 = 32'd78; 
32'd1231: dataIn2 = 32'd96; 
32'd1232: dataIn2 = 32'd31; 
32'd1233: dataIn2 = 32'd41; 
32'd1234: dataIn2 = 32'd44; 
32'd1235: dataIn2 = 32'd1; 
32'd1236: dataIn2 = 32'd47; 
32'd1237: dataIn2 = 32'd98; 
32'd1238: dataIn2 = 32'd4; 
32'd1239: dataIn2 = 32'd21; 
32'd1240: dataIn2 = 32'd60; 
32'd1241: dataIn2 = 32'd57; 
32'd1242: dataIn2 = 32'd8; 
32'd1243: dataIn2 = 32'd40; 
32'd1244: dataIn2 = 32'd36; 
32'd1245: dataIn2 = 32'd52; 
32'd1246: dataIn2 = 32'd72; 
32'd1247: dataIn2 = 32'd99; 
32'd1248: dataIn2 = 32'd46; 
32'd1249: dataIn2 = 32'd84; 
32'd1250: dataIn2 = 32'd14; 
32'd1251: dataIn2 = 32'd12; 
32'd1252: dataIn2 = 32'd61; 
32'd1253: dataIn2 = 32'd42; 
32'd1254: dataIn2 = 32'd51; 
32'd1255: dataIn2 = 32'd62; 
32'd1256: dataIn2 = 32'd86; 
32'd1257: dataIn2 = 32'd2; 
32'd1258: dataIn2 = 32'd5; 
32'd1259: dataIn2 = 32'd17; 
32'd1260: dataIn2 = 32'd81; 
32'd1261: dataIn2 = 32'd96; 
32'd1262: dataIn2 = 32'd18; 
32'd1263: dataIn2 = 32'd25; 
32'd1264: dataIn2 = 32'd97; 
32'd1265: dataIn2 = 32'd10; 
32'd1266: dataIn2 = 32'd82; 
32'd1267: dataIn2 = 32'd35; 
32'd1268: dataIn2 = 32'd27; 
32'd1269: dataIn2 = 32'd96; 
32'd1270: dataIn2 = 32'd96; 
32'd1271: dataIn2 = 32'd79; 
32'd1272: dataIn2 = 32'd46; 
32'd1273: dataIn2 = 32'd15; 
32'd1274: dataIn2 = 32'd44; 
32'd1275: dataIn2 = 32'd13; 
32'd1276: dataIn2 = 32'd23; 
32'd1277: dataIn2 = 32'd35; 
32'd1278: dataIn2 = 32'd47; 
32'd1279: dataIn2 = 32'd28; 
32'd1280: dataIn2 = 32'd61; 
32'd1281: dataIn2 = 32'd95; 
32'd1282: dataIn2 = 32'd71; 
32'd1283: dataIn2 = 32'd95; 
32'd1284: dataIn2 = 32'd71; 
32'd1285: dataIn2 = 32'd17; 
32'd1286: dataIn2 = 32'd40; 
32'd1287: dataIn2 = 32'd16; 
32'd1288: dataIn2 = 32'd61; 
32'd1289: dataIn2 = 32'd52; 
32'd1290: dataIn2 = 32'd39; 
32'd1291: dataIn2 = 32'd77; 
32'd1292: dataIn2 = 32'd52; 
32'd1293: dataIn2 = 32'd36; 
32'd1294: dataIn2 = 32'd72; 
32'd1295: dataIn2 = 32'd9; 
32'd1296: dataIn2 = 32'd68; 
32'd1297: dataIn2 = 32'd24; 
32'd1298: dataIn2 = 32'd26; 
32'd1299: dataIn2 = 32'd20; 
32'd1300: dataIn2 = 32'd45; 
32'd1301: dataIn2 = 32'd31; 
32'd1302: dataIn2 = 32'd87; 
32'd1303: dataIn2 = 32'd20; 
32'd1304: dataIn2 = 32'd67; 
32'd1305: dataIn2 = 32'd10; 
32'd1306: dataIn2 = 32'd6; 
32'd1307: dataIn2 = 32'd33; 
32'd1308: dataIn2 = 32'd22; 
32'd1309: dataIn2 = 32'd8; 
32'd1310: dataIn2 = 32'd33; 
32'd1311: dataIn2 = 32'd59; 
32'd1312: dataIn2 = 32'd92; 
32'd1313: dataIn2 = 32'd77; 
32'd1314: dataIn2 = 32'd39; 
32'd1315: dataIn2 = 32'd46; 
32'd1316: dataIn2 = 32'd23; 
32'd1317: dataIn2 = 32'd79; 
32'd1318: dataIn2 = 32'd31; 
32'd1319: dataIn2 = 32'd28; 
32'd1320: dataIn2 = 32'd7; 
32'd1321: dataIn2 = 32'd46; 
32'd1322: dataIn2 = 32'd24; 
32'd1323: dataIn2 = 32'd89; 
32'd1324: dataIn2 = 32'd17; 
32'd1325: dataIn2 = 32'd57; 
32'd1326: dataIn2 = 32'd85; 
32'd1327: dataIn2 = 32'd15; 
32'd1328: dataIn2 = 32'd64; 
32'd1329: dataIn2 = 32'd74; 
32'd1330: dataIn2 = 32'd30; 
32'd1331: dataIn2 = 32'd17; 
32'd1332: dataIn2 = 32'd25; 
32'd1333: dataIn2 = 32'd30; 
32'd1334: dataIn2 = 32'd97; 
32'd1335: dataIn2 = 32'd48; 
32'd1336: dataIn2 = 32'd52; 
32'd1337: dataIn2 = 32'd58; 
32'd1338: dataIn2 = 32'd10; 
32'd1339: dataIn2 = 32'd57; 
32'd1340: dataIn2 = 32'd13; 
32'd1341: dataIn2 = 32'd82; 
32'd1342: dataIn2 = 32'd47; 
32'd1343: dataIn2 = 32'd61; 
32'd1344: dataIn2 = 32'd68; 
32'd1345: dataIn2 = 32'd36; 
32'd1346: dataIn2 = 32'd29; 
32'd1347: dataIn2 = 32'd0; 
32'd1348: dataIn2 = 32'd74; 
32'd1349: dataIn2 = 32'd88; 
32'd1350: dataIn2 = 32'd78; 
32'd1351: dataIn2 = 32'd35; 
32'd1352: dataIn2 = 32'd60; 
32'd1353: dataIn2 = 32'd93; 
32'd1354: dataIn2 = 32'd21; 
32'd1355: dataIn2 = 32'd22; 
32'd1356: dataIn2 = 32'd2; 
32'd1357: dataIn2 = 32'd4; 
32'd1358: dataIn2 = 32'd32; 
32'd1359: dataIn2 = 32'd54; 
32'd1360: dataIn2 = 32'd52; 
32'd1361: dataIn2 = 32'd81; 
32'd1362: dataIn2 = 32'd80; 
32'd1363: dataIn2 = 32'd19; 
32'd1364: dataIn2 = 32'd48; 
32'd1365: dataIn2 = 32'd72; 
32'd1366: dataIn2 = 32'd67; 
32'd1367: dataIn2 = 32'd24; 
32'd1368: dataIn2 = 32'd8; 
32'd1369: dataIn2 = 32'd50; 
32'd1370: dataIn2 = 32'd66; 
32'd1371: dataIn2 = 32'd16; 
32'd1372: dataIn2 = 32'd21; 
32'd1373: dataIn2 = 32'd83; 
32'd1374: dataIn2 = 32'd78; 
32'd1375: dataIn2 = 32'd7; 
32'd1376: dataIn2 = 32'd23; 
32'd1377: dataIn2 = 32'd63; 
32'd1378: dataIn2 = 32'd2; 
32'd1379: dataIn2 = 32'd2; 
32'd1380: dataIn2 = 32'd10; 
32'd1381: dataIn2 = 32'd27; 
32'd1382: dataIn2 = 32'd45; 
32'd1383: dataIn2 = 32'd33; 
32'd1384: dataIn2 = 32'd43; 
32'd1385: dataIn2 = 32'd32; 
32'd1386: dataIn2 = 32'd96; 
32'd1387: dataIn2 = 32'd12; 
32'd1388: dataIn2 = 32'd20; 
32'd1389: dataIn2 = 32'd19; 
32'd1390: dataIn2 = 32'd10; 
32'd1391: dataIn2 = 32'd53; 
32'd1392: dataIn2 = 32'd99; 
32'd1393: dataIn2 = 32'd96; 
32'd1394: dataIn2 = 32'd90; 
32'd1395: dataIn2 = 32'd46; 
32'd1396: dataIn2 = 32'd46; 
32'd1397: dataIn2 = 32'd71; 
32'd1398: dataIn2 = 32'd87; 
32'd1399: dataIn2 = 32'd5; 
32'd1400: dataIn2 = 32'd39; 
32'd1401: dataIn2 = 32'd50; 
32'd1402: dataIn2 = 32'd70; 
32'd1403: dataIn2 = 32'd78; 
32'd1404: dataIn2 = 32'd34; 
32'd1405: dataIn2 = 32'd88; 
32'd1406: dataIn2 = 32'd57; 
32'd1407: dataIn2 = 32'd17; 
32'd1408: dataIn2 = 32'd18; 
32'd1409: dataIn2 = 32'd28; 
32'd1410: dataIn2 = 32'd39; 
32'd1411: dataIn2 = 32'd27; 
32'd1412: dataIn2 = 32'd97; 
32'd1413: dataIn2 = 32'd72; 
32'd1414: dataIn2 = 32'd43; 
32'd1415: dataIn2 = 32'd45; 
32'd1416: dataIn2 = 32'd67; 
32'd1417: dataIn2 = 32'd25; 
32'd1418: dataIn2 = 32'd10; 
32'd1419: dataIn2 = 32'd49; 
32'd1420: dataIn2 = 32'd10; 
32'd1421: dataIn2 = 32'd43; 
32'd1422: dataIn2 = 32'd76; 
32'd1423: dataIn2 = 32'd97; 
32'd1424: dataIn2 = 32'd12; 
32'd1425: dataIn2 = 32'd7; 
32'd1426: dataIn2 = 32'd9; 
32'd1427: dataIn2 = 32'd58; 
32'd1428: dataIn2 = 32'd57; 
32'd1429: dataIn2 = 32'd60; 
32'd1430: dataIn2 = 32'd42; 
32'd1431: dataIn2 = 32'd62; 
32'd1432: dataIn2 = 32'd9; 
32'd1433: dataIn2 = 32'd29; 
32'd1434: dataIn2 = 32'd72; 
32'd1435: dataIn2 = 32'd19; 
32'd1436: dataIn2 = 32'd20; 
32'd1437: dataIn2 = 32'd1; 
32'd1438: dataIn2 = 32'd4; 
32'd1439: dataIn2 = 32'd42; 
32'd1440: dataIn2 = 32'd86; 
32'd1441: dataIn2 = 32'd73; 
32'd1442: dataIn2 = 32'd97; 
32'd1443: dataIn2 = 32'd53; 
32'd1444: dataIn2 = 32'd32; 
32'd1445: dataIn2 = 32'd33; 
32'd1446: dataIn2 = 32'd18; 
32'd1447: dataIn2 = 32'd58; 
32'd1448: dataIn2 = 32'd99; 
32'd1449: dataIn2 = 32'd34; 
32'd1450: dataIn2 = 32'd59; 
32'd1451: dataIn2 = 32'd91; 
32'd1452: dataIn2 = 32'd31; 
32'd1453: dataIn2 = 32'd0; 
32'd1454: dataIn2 = 32'd93; 
32'd1455: dataIn2 = 32'd81; 
32'd1456: dataIn2 = 32'd35; 
32'd1457: dataIn2 = 32'd35; 
32'd1458: dataIn2 = 32'd68; 
32'd1459: dataIn2 = 32'd74; 
32'd1460: dataIn2 = 32'd98; 
32'd1461: dataIn2 = 32'd67; 
32'd1462: dataIn2 = 32'd31; 
32'd1463: dataIn2 = 32'd54; 
32'd1464: dataIn2 = 32'd7; 
32'd1465: dataIn2 = 32'd8; 
32'd1466: dataIn2 = 32'd67; 
32'd1467: dataIn2 = 32'd93; 
32'd1468: dataIn2 = 32'd37; 
32'd1469: dataIn2 = 32'd56; 
32'd1470: dataIn2 = 32'd55; 
32'd1471: dataIn2 = 32'd89; 
32'd1472: dataIn2 = 32'd3; 
32'd1473: dataIn2 = 32'd74; 
32'd1474: dataIn2 = 32'd21; 
32'd1475: dataIn2 = 32'd5; 
32'd1476: dataIn2 = 32'd36; 
32'd1477: dataIn2 = 32'd99; 
32'd1478: dataIn2 = 32'd19; 
32'd1479: dataIn2 = 32'd100; 
32'd1480: dataIn2 = 32'd20; 
32'd1481: dataIn2 = 32'd63; 
32'd1482: dataIn2 = 32'd73; 
32'd1483: dataIn2 = 32'd73; 
32'd1484: dataIn2 = 32'd10; 
32'd1485: dataIn2 = 32'd41; 
32'd1486: dataIn2 = 32'd90; 
32'd1487: dataIn2 = 32'd62; 
32'd1488: dataIn2 = 32'd50; 
32'd1489: dataIn2 = 32'd14; 
32'd1490: dataIn2 = 32'd4; 
32'd1491: dataIn2 = 32'd30; 
32'd1492: dataIn2 = 32'd26; 
32'd1493: dataIn2 = 32'd94; 
32'd1494: dataIn2 = 32'd66; 
32'd1495: dataIn2 = 32'd63; 
32'd1496: dataIn2 = 32'd12; 
32'd1497: dataIn2 = 32'd60; 
32'd1498: dataIn2 = 32'd67; 
32'd1499: dataIn2 = 32'd5; 
32'd1500: dataIn2 = 32'd73; 
32'd1501: dataIn2 = 32'd93; 
32'd1502: dataIn2 = 32'd28; 
32'd1503: dataIn2 = 32'd31; 
32'd1504: dataIn2 = 32'd90; 
32'd1505: dataIn2 = 32'd29; 
32'd1506: dataIn2 = 32'd15; 
32'd1507: dataIn2 = 32'd10; 
32'd1508: dataIn2 = 32'd62; 
32'd1509: dataIn2 = 32'd34; 
32'd1510: dataIn2 = 32'd51; 
32'd1511: dataIn2 = 32'd69; 
32'd1512: dataIn2 = 32'd88; 
32'd1513: dataIn2 = 32'd31; 
32'd1514: dataIn2 = 32'd99; 
32'd1515: dataIn2 = 32'd32; 
32'd1516: dataIn2 = 32'd25; 
32'd1517: dataIn2 = 32'd59; 
32'd1518: dataIn2 = 32'd0; 
32'd1519: dataIn2 = 32'd87; 
32'd1520: dataIn2 = 32'd62; 
32'd1521: dataIn2 = 32'd31; 
32'd1522: dataIn2 = 32'd63; 
32'd1523: dataIn2 = 32'd81; 
32'd1524: dataIn2 = 32'd49; 
32'd1525: dataIn2 = 32'd52; 
32'd1526: dataIn2 = 32'd8; 
32'd1527: dataIn2 = 32'd30; 
32'd1528: dataIn2 = 32'd52; 
32'd1529: dataIn2 = 32'd78; 
32'd1530: dataIn2 = 32'd94; 
32'd1531: dataIn2 = 32'd62; 
32'd1532: dataIn2 = 32'd8; 
32'd1533: dataIn2 = 32'd97; 
32'd1534: dataIn2 = 32'd52; 
32'd1535: dataIn2 = 32'd35; 
32'd1536: dataIn2 = 32'd74; 
32'd1537: dataIn2 = 32'd55; 
32'd1538: dataIn2 = 32'd21; 
32'd1539: dataIn2 = 32'd94; 
32'd1540: dataIn2 = 32'd56; 
32'd1541: dataIn2 = 32'd13; 
32'd1542: dataIn2 = 32'd54; 
32'd1543: dataIn2 = 32'd87; 
32'd1544: dataIn2 = 32'd75; 
32'd1545: dataIn2 = 32'd84; 
32'd1546: dataIn2 = 32'd35; 
32'd1547: dataIn2 = 32'd1; 
32'd1548: dataIn2 = 32'd8; 
32'd1549: dataIn2 = 32'd40; 
32'd1550: dataIn2 = 32'd47; 
32'd1551: dataIn2 = 32'd94; 
32'd1552: dataIn2 = 32'd47; 
32'd1553: dataIn2 = 32'd72; 
32'd1554: dataIn2 = 32'd1; 
32'd1555: dataIn2 = 32'd32; 
32'd1556: dataIn2 = 32'd12; 
32'd1557: dataIn2 = 32'd19; 
32'd1558: dataIn2 = 32'd65; 
32'd1559: dataIn2 = 32'd30; 
32'd1560: dataIn2 = 32'd54; 
32'd1561: dataIn2 = 32'd95; 
32'd1562: dataIn2 = 32'd48; 
32'd1563: dataIn2 = 32'd48; 
32'd1564: dataIn2 = 32'd79; 
32'd1565: dataIn2 = 32'd76; 
32'd1566: dataIn2 = 32'd64; 
32'd1567: dataIn2 = 32'd75; 
32'd1568: dataIn2 = 32'd33; 
32'd1569: dataIn2 = 32'd35; 
32'd1570: dataIn2 = 32'd8; 
32'd1571: dataIn2 = 32'd22; 
32'd1572: dataIn2 = 32'd16; 
32'd1573: dataIn2 = 32'd65; 
32'd1574: dataIn2 = 32'd70; 
32'd1575: dataIn2 = 32'd22; 
32'd1576: dataIn2 = 32'd61; 
32'd1577: dataIn2 = 32'd32; 
32'd1578: dataIn2 = 32'd93; 
32'd1579: dataIn2 = 32'd14; 
32'd1580: dataIn2 = 32'd21; 
32'd1581: dataIn2 = 32'd72; 
32'd1582: dataIn2 = 32'd34; 
32'd1583: dataIn2 = 32'd1; 
32'd1584: dataIn2 = 32'd69; 
32'd1585: dataIn2 = 32'd3; 
32'd1586: dataIn2 = 32'd29; 
32'd1587: dataIn2 = 32'd53; 
32'd1588: dataIn2 = 32'd21; 
32'd1589: dataIn2 = 32'd96; 
32'd1590: dataIn2 = 32'd13; 
32'd1591: dataIn2 = 32'd73; 
32'd1592: dataIn2 = 32'd70; 
32'd1593: dataIn2 = 32'd76; 
32'd1594: dataIn2 = 32'd60; 
32'd1595: dataIn2 = 32'd63; 
32'd1596: dataIn2 = 32'd58; 
32'd1597: dataIn2 = 32'd17; 
32'd1598: dataIn2 = 32'd12; 
32'd1599: dataIn2 = 32'd10; 
32'd1600: dataIn2 = 32'd47; 
32'd1601: dataIn2 = 32'd66; 
32'd1602: dataIn2 = 32'd90; 
32'd1603: dataIn2 = 32'd42; 
32'd1604: dataIn2 = 32'd84; 
32'd1605: dataIn2 = 32'd36; 
32'd1606: dataIn2 = 32'd90; 
32'd1607: dataIn2 = 32'd52; 
32'd1608: dataIn2 = 32'd16; 
32'd1609: dataIn2 = 32'd2; 
32'd1610: dataIn2 = 32'd75; 
32'd1611: dataIn2 = 32'd12; 
32'd1612: dataIn2 = 32'd37; 
32'd1613: dataIn2 = 32'd70; 
32'd1614: dataIn2 = 32'd45; 
32'd1615: dataIn2 = 32'd4; 
32'd1616: dataIn2 = 32'd19; 
32'd1617: dataIn2 = 32'd100; 
32'd1618: dataIn2 = 32'd69; 
32'd1619: dataIn2 = 32'd63; 
32'd1620: dataIn2 = 32'd87; 
32'd1621: dataIn2 = 32'd45; 
32'd1622: dataIn2 = 32'd80; 
32'd1623: dataIn2 = 32'd3; 
32'd1624: dataIn2 = 32'd37; 
32'd1625: dataIn2 = 32'd81; 
32'd1626: dataIn2 = 32'd69; 
32'd1627: dataIn2 = 32'd55; 
32'd1628: dataIn2 = 32'd48; 
32'd1629: dataIn2 = 32'd8; 
32'd1630: dataIn2 = 32'd9; 
32'd1631: dataIn2 = 32'd69; 
32'd1632: dataIn2 = 32'd96; 
32'd1633: dataIn2 = 32'd59; 
32'd1634: dataIn2 = 32'd18; 
32'd1635: dataIn2 = 32'd28; 
32'd1636: dataIn2 = 32'd85; 
32'd1637: dataIn2 = 32'd67; 
32'd1638: dataIn2 = 32'd81; 
32'd1639: dataIn2 = 32'd41; 
32'd1640: dataIn2 = 32'd24; 
32'd1641: dataIn2 = 32'd30; 
32'd1642: dataIn2 = 32'd80; 
32'd1643: dataIn2 = 32'd16; 
32'd1644: dataIn2 = 32'd98; 
32'd1645: dataIn2 = 32'd80; 
32'd1646: dataIn2 = 32'd93; 
32'd1647: dataIn2 = 32'd56; 
32'd1648: dataIn2 = 32'd42; 
32'd1649: dataIn2 = 32'd48; 
32'd1650: dataIn2 = 32'd96; 
32'd1651: dataIn2 = 32'd61; 
32'd1652: dataIn2 = 32'd26; 
32'd1653: dataIn2 = 32'd20; 
32'd1654: dataIn2 = 32'd12; 
32'd1655: dataIn2 = 32'd18; 
32'd1656: dataIn2 = 32'd14; 
32'd1657: dataIn2 = 32'd58; 
32'd1658: dataIn2 = 32'd46; 
32'd1659: dataIn2 = 32'd15; 
32'd1660: dataIn2 = 32'd16; 
32'd1661: dataIn2 = 32'd35; 
32'd1662: dataIn2 = 32'd77; 
32'd1663: dataIn2 = 32'd18; 
32'd1664: dataIn2 = 32'd96; 
32'd1665: dataIn2 = 32'd26; 
32'd1666: dataIn2 = 32'd73; 
32'd1667: dataIn2 = 32'd31; 
32'd1668: dataIn2 = 32'd67; 
32'd1669: dataIn2 = 32'd9; 
32'd1670: dataIn2 = 32'd92; 
32'd1671: dataIn2 = 32'd78; 
32'd1672: dataIn2 = 32'd86; 
32'd1673: dataIn2 = 32'd22; 
32'd1674: dataIn2 = 32'd97; 
32'd1675: dataIn2 = 32'd69; 
32'd1676: dataIn2 = 32'd68; 
32'd1677: dataIn2 = 32'd9; 
32'd1678: dataIn2 = 32'd9; 
32'd1679: dataIn2 = 32'd80; 
32'd1680: dataIn2 = 32'd47; 
32'd1681: dataIn2 = 32'd2; 
32'd1682: dataIn2 = 32'd87; 
32'd1683: dataIn2 = 32'd60; 
32'd1684: dataIn2 = 32'd27; 
32'd1685: dataIn2 = 32'd35; 
32'd1686: dataIn2 = 32'd85; 
32'd1687: dataIn2 = 32'd4; 
32'd1688: dataIn2 = 32'd97; 
32'd1689: dataIn2 = 32'd47; 
32'd1690: dataIn2 = 32'd69; 
32'd1691: dataIn2 = 32'd26; 
32'd1692: dataIn2 = 32'd94; 
32'd1693: dataIn2 = 32'd4; 
32'd1694: dataIn2 = 32'd91; 
32'd1695: dataIn2 = 32'd32; 
32'd1696: dataIn2 = 32'd16; 
32'd1697: dataIn2 = 32'd63; 
32'd1698: dataIn2 = 32'd98; 
32'd1699: dataIn2 = 32'd28; 
32'd1700: dataIn2 = 32'd17; 
32'd1701: dataIn2 = 32'd29; 
32'd1702: dataIn2 = 32'd25; 
32'd1703: dataIn2 = 32'd6; 
32'd1704: dataIn2 = 32'd27; 
32'd1705: dataIn2 = 32'd75; 
32'd1706: dataIn2 = 32'd100; 
32'd1707: dataIn2 = 32'd73; 
32'd1708: dataIn2 = 32'd51; 
32'd1709: dataIn2 = 32'd2; 
32'd1710: dataIn2 = 32'd41; 
32'd1711: dataIn2 = 32'd36; 
32'd1712: dataIn2 = 32'd45; 
32'd1713: dataIn2 = 32'd68; 
32'd1714: dataIn2 = 32'd21; 
32'd1715: dataIn2 = 32'd82; 
32'd1716: dataIn2 = 32'd30; 
32'd1717: dataIn2 = 32'd90; 
32'd1718: dataIn2 = 32'd24; 
32'd1719: dataIn2 = 32'd3; 
32'd1720: dataIn2 = 32'd41; 
32'd1721: dataIn2 = 32'd71; 
32'd1722: dataIn2 = 32'd73; 
32'd1723: dataIn2 = 32'd39; 
32'd1724: dataIn2 = 32'd91; 
32'd1725: dataIn2 = 32'd97; 
32'd1726: dataIn2 = 32'd0; 
32'd1727: dataIn2 = 32'd21; 
32'd1728: dataIn2 = 32'd25; 
32'd1729: dataIn2 = 32'd9; 
32'd1730: dataIn2 = 32'd99; 
32'd1731: dataIn2 = 32'd99; 
32'd1732: dataIn2 = 32'd11; 
32'd1733: dataIn2 = 32'd63; 
32'd1734: dataIn2 = 32'd49; 
32'd1735: dataIn2 = 32'd57; 
32'd1736: dataIn2 = 32'd3; 
32'd1737: dataIn2 = 32'd75; 
32'd1738: dataIn2 = 32'd72; 
32'd1739: dataIn2 = 32'd49; 
32'd1740: dataIn2 = 32'd42; 
32'd1741: dataIn2 = 32'd26; 
32'd1742: dataIn2 = 32'd27; 
32'd1743: dataIn2 = 32'd77; 
32'd1744: dataIn2 = 32'd30; 
32'd1745: dataIn2 = 32'd62; 
32'd1746: dataIn2 = 32'd99; 
32'd1747: dataIn2 = 32'd0; 
32'd1748: dataIn2 = 32'd53; 
32'd1749: dataIn2 = 32'd90; 
32'd1750: dataIn2 = 32'd5; 
32'd1751: dataIn2 = 32'd11; 
32'd1752: dataIn2 = 32'd58; 
32'd1753: dataIn2 = 32'd96; 
32'd1754: dataIn2 = 32'd50; 
32'd1755: dataIn2 = 32'd54; 
32'd1756: dataIn2 = 32'd45; 
32'd1757: dataIn2 = 32'd88; 
32'd1758: dataIn2 = 32'd93; 
32'd1759: dataIn2 = 32'd44; 
32'd1760: dataIn2 = 32'd93; 
32'd1761: dataIn2 = 32'd39; 
32'd1762: dataIn2 = 32'd91; 
32'd1763: dataIn2 = 32'd7; 
32'd1764: dataIn2 = 32'd24; 
32'd1765: dataIn2 = 32'd29; 
32'd1766: dataIn2 = 32'd53; 
32'd1767: dataIn2 = 32'd14; 
32'd1768: dataIn2 = 32'd58; 
32'd1769: dataIn2 = 32'd14; 
32'd1770: dataIn2 = 32'd2; 
32'd1771: dataIn2 = 32'd96; 
32'd1772: dataIn2 = 32'd43; 
32'd1773: dataIn2 = 32'd42; 
32'd1774: dataIn2 = 32'd47; 
32'd1775: dataIn2 = 32'd66; 
32'd1776: dataIn2 = 32'd6; 
32'd1777: dataIn2 = 32'd85; 
32'd1778: dataIn2 = 32'd34; 
32'd1779: dataIn2 = 32'd24; 
32'd1780: dataIn2 = 32'd74; 
32'd1781: dataIn2 = 32'd1; 
32'd1782: dataIn2 = 32'd14; 
32'd1783: dataIn2 = 32'd58; 
32'd1784: dataIn2 = 32'd95; 
32'd1785: dataIn2 = 32'd76; 
32'd1786: dataIn2 = 32'd82; 
32'd1787: dataIn2 = 32'd15; 
32'd1788: dataIn2 = 32'd53; 
32'd1789: dataIn2 = 32'd44; 
32'd1790: dataIn2 = 32'd87; 
32'd1791: dataIn2 = 32'd77; 
32'd1792: dataIn2 = 32'd55; 
32'd1793: dataIn2 = 32'd68; 
32'd1794: dataIn2 = 32'd23; 
32'd1795: dataIn2 = 32'd33; 
32'd1796: dataIn2 = 32'd23; 
32'd1797: dataIn2 = 32'd87; 
32'd1798: dataIn2 = 32'd55; 
32'd1799: dataIn2 = 32'd44; 
32'd1800: dataIn2 = 32'd40; 
32'd1801: dataIn2 = 32'd52; 
32'd1802: dataIn2 = 32'd58; 
32'd1803: dataIn2 = 32'd15; 
32'd1804: dataIn2 = 32'd46; 
32'd1805: dataIn2 = 32'd79; 
32'd1806: dataIn2 = 32'd96; 
32'd1807: dataIn2 = 32'd76; 
32'd1808: dataIn2 = 32'd42; 
32'd1809: dataIn2 = 32'd54; 
32'd1810: dataIn2 = 32'd78; 
32'd1811: dataIn2 = 32'd33; 
32'd1812: dataIn2 = 32'd60; 
32'd1813: dataIn2 = 32'd19; 
32'd1814: dataIn2 = 32'd25; 
32'd1815: dataIn2 = 32'd62; 
32'd1816: dataIn2 = 32'd2; 
32'd1817: dataIn2 = 32'd19; 
32'd1818: dataIn2 = 32'd49; 
32'd1819: dataIn2 = 32'd27; 
32'd1820: dataIn2 = 32'd59; 
32'd1821: dataIn2 = 32'd54; 
32'd1822: dataIn2 = 32'd26; 
32'd1823: dataIn2 = 32'd19; 
32'd1824: dataIn2 = 32'd24; 
32'd1825: dataIn2 = 32'd30; 
32'd1826: dataIn2 = 32'd83; 
32'd1827: dataIn2 = 32'd71; 
32'd1828: dataIn2 = 32'd55; 
32'd1829: dataIn2 = 32'd31; 
32'd1830: dataIn2 = 32'd57; 
32'd1831: dataIn2 = 32'd65; 
32'd1832: dataIn2 = 32'd2; 
32'd1833: dataIn2 = 32'd54; 
32'd1834: dataIn2 = 32'd31; 
32'd1835: dataIn2 = 32'd1; 
32'd1836: dataIn2 = 32'd14; 
32'd1837: dataIn2 = 32'd10; 
32'd1838: dataIn2 = 32'd21; 
32'd1839: dataIn2 = 32'd62; 
32'd1840: dataIn2 = 32'd28; 
32'd1841: dataIn2 = 32'd86; 
32'd1842: dataIn2 = 32'd81; 
32'd1843: dataIn2 = 32'd95; 
32'd1844: dataIn2 = 32'd8; 
32'd1845: dataIn2 = 32'd45; 
32'd1846: dataIn2 = 32'd7; 
32'd1847: dataIn2 = 32'd14; 
32'd1848: dataIn2 = 32'd16; 
32'd1849: dataIn2 = 32'd85; 
32'd1850: dataIn2 = 32'd91; 
32'd1851: dataIn2 = 32'd6; 
32'd1852: dataIn2 = 32'd56; 
32'd1853: dataIn2 = 32'd59; 
32'd1854: dataIn2 = 32'd76; 
32'd1855: dataIn2 = 32'd41; 
32'd1856: dataIn2 = 32'd90; 
32'd1857: dataIn2 = 32'd65; 
32'd1858: dataIn2 = 32'd86; 
32'd1859: dataIn2 = 32'd58; 
32'd1860: dataIn2 = 32'd44; 
32'd1861: dataIn2 = 32'd48; 
32'd1862: dataIn2 = 32'd4; 
32'd1863: dataIn2 = 32'd19; 
32'd1864: dataIn2 = 32'd81; 
32'd1865: dataIn2 = 32'd63; 
32'd1866: dataIn2 = 32'd68; 
32'd1867: dataIn2 = 32'd98; 
32'd1868: dataIn2 = 32'd54; 
32'd1869: dataIn2 = 32'd98; 
32'd1870: dataIn2 = 32'd90; 
32'd1871: dataIn2 = 32'd8; 
32'd1872: dataIn2 = 32'd59; 
32'd1873: dataIn2 = 32'd4; 
32'd1874: dataIn2 = 32'd59; 
32'd1875: dataIn2 = 32'd76; 
32'd1876: dataIn2 = 32'd77; 
32'd1877: dataIn2 = 32'd91; 
32'd1878: dataIn2 = 32'd34; 
32'd1879: dataIn2 = 32'd30; 
32'd1880: dataIn2 = 32'd46; 
32'd1881: dataIn2 = 32'd27; 
32'd1882: dataIn2 = 32'd6; 
32'd1883: dataIn2 = 32'd25; 
32'd1884: dataIn2 = 32'd62; 
32'd1885: dataIn2 = 32'd41; 
32'd1886: dataIn2 = 32'd16; 
32'd1887: dataIn2 = 32'd100; 
32'd1888: dataIn2 = 32'd35; 
32'd1889: dataIn2 = 32'd91; 
32'd1890: dataIn2 = 32'd94; 
32'd1891: dataIn2 = 32'd37; 
32'd1892: dataIn2 = 32'd74; 
32'd1893: dataIn2 = 32'd79; 
32'd1894: dataIn2 = 32'd95; 
32'd1895: dataIn2 = 32'd62; 
32'd1896: dataIn2 = 32'd7; 
32'd1897: dataIn2 = 32'd67; 
32'd1898: dataIn2 = 32'd81; 
32'd1899: dataIn2 = 32'd65; 
32'd1900: dataIn2 = 32'd94; 
32'd1901: dataIn2 = 32'd12; 
32'd1902: dataIn2 = 32'd5; 
32'd1903: dataIn2 = 32'd89; 
32'd1904: dataIn2 = 32'd47; 
32'd1905: dataIn2 = 32'd42; 
32'd1906: dataIn2 = 32'd78; 
32'd1907: dataIn2 = 32'd99; 
32'd1908: dataIn2 = 32'd18; 
32'd1909: dataIn2 = 32'd37; 
32'd1910: dataIn2 = 32'd91; 
32'd1911: dataIn2 = 32'd5; 
32'd1912: dataIn2 = 32'd6; 
32'd1913: dataIn2 = 32'd78; 
32'd1914: dataIn2 = 32'd17; 
32'd1915: dataIn2 = 32'd10; 
32'd1916: dataIn2 = 32'd83; 
32'd1917: dataIn2 = 32'd4; 
32'd1918: dataIn2 = 32'd71; 
32'd1919: dataIn2 = 32'd26; 
32'd1920: dataIn2 = 32'd92; 
32'd1921: dataIn2 = 32'd99; 
32'd1922: dataIn2 = 32'd40; 
32'd1923: dataIn2 = 32'd57; 
32'd1924: dataIn2 = 32'd92; 
32'd1925: dataIn2 = 32'd78; 
32'd1926: dataIn2 = 32'd43; 
32'd1927: dataIn2 = 32'd86; 
32'd1928: dataIn2 = 32'd32; 
32'd1929: dataIn2 = 32'd29; 
32'd1930: dataIn2 = 32'd30; 
32'd1931: dataIn2 = 32'd38; 
32'd1932: dataIn2 = 32'd60; 
32'd1933: dataIn2 = 32'd60; 
32'd1934: dataIn2 = 32'd56; 
32'd1935: dataIn2 = 32'd5; 
32'd1936: dataIn2 = 32'd43; 
32'd1937: dataIn2 = 32'd43; 
32'd1938: dataIn2 = 32'd76; 
32'd1939: dataIn2 = 32'd63; 
32'd1940: dataIn2 = 32'd12; 
32'd1941: dataIn2 = 32'd30; 
32'd1942: dataIn2 = 32'd35; 
32'd1943: dataIn2 = 32'd87; 
32'd1944: dataIn2 = 32'd74; 
32'd1945: dataIn2 = 32'd54; 
32'd1946: dataIn2 = 32'd89; 
32'd1947: dataIn2 = 32'd23; 
32'd1948: dataIn2 = 32'd51; 
32'd1949: dataIn2 = 32'd95; 
32'd1950: dataIn2 = 32'd31; 
32'd1951: dataIn2 = 32'd23; 
32'd1952: dataIn2 = 32'd31; 
32'd1953: dataIn2 = 32'd32; 
32'd1954: dataIn2 = 32'd31; 
32'd1955: dataIn2 = 32'd99; 
32'd1956: dataIn2 = 32'd87; 
32'd1957: dataIn2 = 32'd49; 
32'd1958: dataIn2 = 32'd50; 
32'd1959: dataIn2 = 32'd11; 
32'd1960: dataIn2 = 32'd59; 
32'd1961: dataIn2 = 32'd68; 
32'd1962: dataIn2 = 32'd39; 
32'd1963: dataIn2 = 32'd11; 
32'd1964: dataIn2 = 32'd90; 
32'd1965: dataIn2 = 32'd45; 
32'd1966: dataIn2 = 32'd13; 
32'd1967: dataIn2 = 32'd83; 
32'd1968: dataIn2 = 32'd32; 
32'd1969: dataIn2 = 32'd94; 
32'd1970: dataIn2 = 32'd51; 
32'd1971: dataIn2 = 32'd71; 
32'd1972: dataIn2 = 32'd86; 
32'd1973: dataIn2 = 32'd83; 
32'd1974: dataIn2 = 32'd56; 
32'd1975: dataIn2 = 32'd68; 
32'd1976: dataIn2 = 32'd50; 
32'd1977: dataIn2 = 32'd36; 
32'd1978: dataIn2 = 32'd50; 
32'd1979: dataIn2 = 32'd37; 
32'd1980: dataIn2 = 32'd62; 
32'd1981: dataIn2 = 32'd1; 
32'd1982: dataIn2 = 32'd8; 
32'd1983: dataIn2 = 32'd99; 
32'd1984: dataIn2 = 32'd72; 
32'd1985: dataIn2 = 32'd55; 
32'd1986: dataIn2 = 32'd12; 
32'd1987: dataIn2 = 32'd56; 
32'd1988: dataIn2 = 32'd50; 
32'd1989: dataIn2 = 32'd82; 
32'd1990: dataIn2 = 32'd85; 
32'd1991: dataIn2 = 32'd30; 
32'd1992: dataIn2 = 32'd93; 
32'd1993: dataIn2 = 32'd7; 
32'd1994: dataIn2 = 32'd29; 
32'd1995: dataIn2 = 32'd71; 
32'd1996: dataIn2 = 32'd37; 
32'd1997: dataIn2 = 32'd6; 
32'd1998: dataIn2 = 32'd22; 
32'd1999: dataIn2 = 32'd19; 
32'd2000: dataIn2 = 32'd10; 
32'd2001: dataIn2 = 32'd16; 
32'd2002: dataIn2 = 32'd3; 
32'd2003: dataIn2 = 32'd37; 
32'd2004: dataIn2 = 32'd12; 
32'd2005: dataIn2 = 32'd79; 
32'd2006: dataIn2 = 32'd27; 
32'd2007: dataIn2 = 32'd50; 
32'd2008: dataIn2 = 32'd69; 
32'd2009: dataIn2 = 32'd67; 
32'd2010: dataIn2 = 32'd82; 
32'd2011: dataIn2 = 32'd100; 
32'd2012: dataIn2 = 32'd75; 
32'd2013: dataIn2 = 32'd22; 
32'd2014: dataIn2 = 32'd14; 
32'd2015: dataIn2 = 32'd56; 
32'd2016: dataIn2 = 32'd91; 
32'd2017: dataIn2 = 32'd48; 
32'd2018: dataIn2 = 32'd100; 
32'd2019: dataIn2 = 32'd100; 
32'd2020: dataIn2 = 32'd26; 
32'd2021: dataIn2 = 32'd11; 
32'd2022: dataIn2 = 32'd76; 
32'd2023: dataIn2 = 32'd60; 
32'd2024: dataIn2 = 32'd71; 
32'd2025: dataIn2 = 32'd8; 
32'd2026: dataIn2 = 32'd86; 
32'd2027: dataIn2 = 32'd35; 
32'd2028: dataIn2 = 32'd24; 
32'd2029: dataIn2 = 32'd12; 
32'd2030: dataIn2 = 32'd36; 
32'd2031: dataIn2 = 32'd4; 
32'd2032: dataIn2 = 32'd21; 
32'd2033: dataIn2 = 32'd48; 
32'd2034: dataIn2 = 32'd65; 
32'd2035: dataIn2 = 32'd99; 
32'd2036: dataIn2 = 32'd44; 
32'd2037: dataIn2 = 32'd42; 
32'd2038: dataIn2 = 32'd54; 
32'd2039: dataIn2 = 32'd45; 
32'd2040: dataIn2 = 32'd100; 
32'd2041: dataIn2 = 32'd97; 
32'd2042: dataIn2 = 32'd9; 
32'd2043: dataIn2 = 32'd7; 
32'd2044: dataIn2 = 32'd0; 
32'd2045: dataIn2 = 32'd32; 
32'd2046: dataIn2 = 32'd70; 
32'd2047: dataIn2 = 32'd5; 
32'd2048: dataIn2 = 32'd52; 
32'd2049: dataIn2 = 32'd34; 
32'd2050: dataIn2 = 32'd11; 
32'd2051: dataIn2 = 32'd5; 
32'd2052: dataIn2 = 32'd31; 
32'd2053: dataIn2 = 32'd24; 
32'd2054: dataIn2 = 32'd21; 
32'd2055: dataIn2 = 32'd35; 
32'd2056: dataIn2 = 32'd66; 
32'd2057: dataIn2 = 32'd7; 
32'd2058: dataIn2 = 32'd86; 
32'd2059: dataIn2 = 32'd25; 
32'd2060: dataIn2 = 32'd63; 
32'd2061: dataIn2 = 32'd70; 
32'd2062: dataIn2 = 32'd85; 
32'd2063: dataIn2 = 32'd1; 
32'd2064: dataIn2 = 32'd52; 
32'd2065: dataIn2 = 32'd23; 
32'd2066: dataIn2 = 32'd87; 
32'd2067: dataIn2 = 32'd5; 
32'd2068: dataIn2 = 32'd84; 
32'd2069: dataIn2 = 32'd40; 
32'd2070: dataIn2 = 32'd45; 
32'd2071: dataIn2 = 32'd54; 
32'd2072: dataIn2 = 32'd85; 
32'd2073: dataIn2 = 32'd93; 
32'd2074: dataIn2 = 32'd100; 
32'd2075: dataIn2 = 32'd63; 
32'd2076: dataIn2 = 32'd52; 
32'd2077: dataIn2 = 32'd56; 
32'd2078: dataIn2 = 32'd22; 
32'd2079: dataIn2 = 32'd90; 
32'd2080: dataIn2 = 32'd27; 
32'd2081: dataIn2 = 32'd16; 
32'd2082: dataIn2 = 32'd93; 
32'd2083: dataIn2 = 32'd77; 
32'd2084: dataIn2 = 32'd97; 
32'd2085: dataIn2 = 32'd50; 
32'd2086: dataIn2 = 32'd19; 
32'd2087: dataIn2 = 32'd17; 
32'd2088: dataIn2 = 32'd79; 
32'd2089: dataIn2 = 32'd77; 
32'd2090: dataIn2 = 32'd24; 
32'd2091: dataIn2 = 32'd28; 
32'd2092: dataIn2 = 32'd37; 
32'd2093: dataIn2 = 32'd29; 
32'd2094: dataIn2 = 32'd29; 
32'd2095: dataIn2 = 32'd37; 
32'd2096: dataIn2 = 32'd61; 
32'd2097: dataIn2 = 32'd54; 
32'd2098: dataIn2 = 32'd28; 
32'd2099: dataIn2 = 32'd53; 
32'd2100: dataIn2 = 32'd94; 
32'd2101: dataIn2 = 32'd70; 
32'd2102: dataIn2 = 32'd66; 
32'd2103: dataIn2 = 32'd15; 
32'd2104: dataIn2 = 32'd1; 
32'd2105: dataIn2 = 32'd53; 
32'd2106: dataIn2 = 32'd5; 
32'd2107: dataIn2 = 32'd41; 
32'd2108: dataIn2 = 32'd17; 
32'd2109: dataIn2 = 32'd98; 
32'd2110: dataIn2 = 32'd87; 
32'd2111: dataIn2 = 32'd29; 
32'd2112: dataIn2 = 32'd61; 
32'd2113: dataIn2 = 32'd97; 
32'd2114: dataIn2 = 32'd96; 
32'd2115: dataIn2 = 32'd19; 
32'd2116: dataIn2 = 32'd27; 
32'd2117: dataIn2 = 32'd80; 
32'd2118: dataIn2 = 32'd1; 
32'd2119: dataIn2 = 32'd21; 
32'd2120: dataIn2 = 32'd37; 
32'd2121: dataIn2 = 32'd31; 
32'd2122: dataIn2 = 32'd57; 
32'd2123: dataIn2 = 32'd46; 
32'd2124: dataIn2 = 32'd6; 
32'd2125: dataIn2 = 32'd10; 
32'd2126: dataIn2 = 32'd50; 
32'd2127: dataIn2 = 32'd58; 
32'd2128: dataIn2 = 32'd66; 
32'd2129: dataIn2 = 32'd34; 
32'd2130: dataIn2 = 32'd73; 
32'd2131: dataIn2 = 32'd1; 
32'd2132: dataIn2 = 32'd36; 
32'd2133: dataIn2 = 32'd24; 
32'd2134: dataIn2 = 32'd11; 
32'd2135: dataIn2 = 32'd6; 
32'd2136: dataIn2 = 32'd11; 
32'd2137: dataIn2 = 32'd27; 
32'd2138: dataIn2 = 32'd40; 
32'd2139: dataIn2 = 32'd27; 
32'd2140: dataIn2 = 32'd61; 
32'd2141: dataIn2 = 32'd63; 
32'd2142: dataIn2 = 32'd73; 
32'd2143: dataIn2 = 32'd21; 
32'd2144: dataIn2 = 32'd63; 
32'd2145: dataIn2 = 32'd22; 
32'd2146: dataIn2 = 32'd82; 
32'd2147: dataIn2 = 32'd90; 
32'd2148: dataIn2 = 32'd92; 
32'd2149: dataIn2 = 32'd55; 
32'd2150: dataIn2 = 32'd92; 
32'd2151: dataIn2 = 32'd25; 
32'd2152: dataIn2 = 32'd16; 
32'd2153: dataIn2 = 32'd15; 
32'd2154: dataIn2 = 32'd32; 
32'd2155: dataIn2 = 32'd96; 
32'd2156: dataIn2 = 32'd71; 
32'd2157: dataIn2 = 32'd82; 
32'd2158: dataIn2 = 32'd70; 
32'd2159: dataIn2 = 32'd43; 
32'd2160: dataIn2 = 32'd67; 
32'd2161: dataIn2 = 32'd30; 
32'd2162: dataIn2 = 32'd96; 
32'd2163: dataIn2 = 32'd31; 
32'd2164: dataIn2 = 32'd81; 
32'd2165: dataIn2 = 32'd12; 
32'd2166: dataIn2 = 32'd92; 
32'd2167: dataIn2 = 32'd45; 
32'd2168: dataIn2 = 32'd86; 
32'd2169: dataIn2 = 32'd52; 
32'd2170: dataIn2 = 32'd96; 
32'd2171: dataIn2 = 32'd18; 
32'd2172: dataIn2 = 32'd29; 
32'd2173: dataIn2 = 32'd69; 
32'd2174: dataIn2 = 32'd93; 
32'd2175: dataIn2 = 32'd84; 
32'd2176: dataIn2 = 32'd93; 
32'd2177: dataIn2 = 32'd11; 
32'd2178: dataIn2 = 32'd36; 
32'd2179: dataIn2 = 32'd91; 
32'd2180: dataIn2 = 32'd34; 
32'd2181: dataIn2 = 32'd44; 
32'd2182: dataIn2 = 32'd53; 
32'd2183: dataIn2 = 32'd89; 
32'd2184: dataIn2 = 32'd58; 
32'd2185: dataIn2 = 32'd40; 
32'd2186: dataIn2 = 32'd70; 
32'd2187: dataIn2 = 32'd92; 
32'd2188: dataIn2 = 32'd91; 
32'd2189: dataIn2 = 32'd32; 
32'd2190: dataIn2 = 32'd60; 
32'd2191: dataIn2 = 32'd84; 
32'd2192: dataIn2 = 32'd44; 
32'd2193: dataIn2 = 32'd84; 
32'd2194: dataIn2 = 32'd40; 
32'd2195: dataIn2 = 32'd28; 
32'd2196: dataIn2 = 32'd77; 
32'd2197: dataIn2 = 32'd48; 
32'd2198: dataIn2 = 32'd74; 
32'd2199: dataIn2 = 32'd24; 
32'd2200: dataIn2 = 32'd89; 
32'd2201: dataIn2 = 32'd36; 
32'd2202: dataIn2 = 32'd29; 
32'd2203: dataIn2 = 32'd36; 
32'd2204: dataIn2 = 32'd52; 
32'd2205: dataIn2 = 32'd88; 
32'd2206: dataIn2 = 32'd64; 
32'd2207: dataIn2 = 32'd39; 
32'd2208: dataIn2 = 32'd66; 
32'd2209: dataIn2 = 32'd74; 
32'd2210: dataIn2 = 32'd0; 
32'd2211: dataIn2 = 32'd65; 
32'd2212: dataIn2 = 32'd25; 
32'd2213: dataIn2 = 32'd21; 
32'd2214: dataIn2 = 32'd38; 
32'd2215: dataIn2 = 32'd20; 
32'd2216: dataIn2 = 32'd76; 
32'd2217: dataIn2 = 32'd93; 
32'd2218: dataIn2 = 32'd50; 
32'd2219: dataIn2 = 32'd79; 
32'd2220: dataIn2 = 32'd26; 
32'd2221: dataIn2 = 32'd26; 
32'd2222: dataIn2 = 32'd4; 
32'd2223: dataIn2 = 32'd45; 
32'd2224: dataIn2 = 32'd22; 
32'd2225: dataIn2 = 32'd97; 
32'd2226: dataIn2 = 32'd9; 
32'd2227: dataIn2 = 32'd53; 
32'd2228: dataIn2 = 32'd53; 
32'd2229: dataIn2 = 32'd53; 
32'd2230: dataIn2 = 32'd59; 
32'd2231: dataIn2 = 32'd74; 
32'd2232: dataIn2 = 32'd52; 
32'd2233: dataIn2 = 32'd59; 
32'd2234: dataIn2 = 32'd42; 
32'd2235: dataIn2 = 32'd7; 
32'd2236: dataIn2 = 32'd2; 
32'd2237: dataIn2 = 32'd86; 
32'd2238: dataIn2 = 32'd91; 
32'd2239: dataIn2 = 32'd30; 
32'd2240: dataIn2 = 32'd89; 
32'd2241: dataIn2 = 32'd67; 
32'd2242: dataIn2 = 32'd22; 
32'd2243: dataIn2 = 32'd59; 
32'd2244: dataIn2 = 32'd0; 
32'd2245: dataIn2 = 32'd70; 
32'd2246: dataIn2 = 32'd3; 
32'd2247: dataIn2 = 32'd58; 
32'd2248: dataIn2 = 32'd47; 
32'd2249: dataIn2 = 32'd59; 
32'd2250: dataIn2 = 32'd18; 
32'd2251: dataIn2 = 32'd43; 
32'd2252: dataIn2 = 32'd25; 
32'd2253: dataIn2 = 32'd23; 
32'd2254: dataIn2 = 32'd22; 
32'd2255: dataIn2 = 32'd68; 
32'd2256: dataIn2 = 32'd30; 
32'd2257: dataIn2 = 32'd45; 
32'd2258: dataIn2 = 32'd34; 
32'd2259: dataIn2 = 32'd7; 
32'd2260: dataIn2 = 32'd40; 
32'd2261: dataIn2 = 32'd92; 
32'd2262: dataIn2 = 32'd64; 
32'd2263: dataIn2 = 32'd58; 
32'd2264: dataIn2 = 32'd62; 
32'd2265: dataIn2 = 32'd56; 
32'd2266: dataIn2 = 32'd79; 
32'd2267: dataIn2 = 32'd61; 
32'd2268: dataIn2 = 32'd62; 
32'd2269: dataIn2 = 32'd66; 
32'd2270: dataIn2 = 32'd50; 
32'd2271: dataIn2 = 32'd60; 
32'd2272: dataIn2 = 32'd47; 
32'd2273: dataIn2 = 32'd99; 
32'd2274: dataIn2 = 32'd94; 
32'd2275: dataIn2 = 32'd45; 
32'd2276: dataIn2 = 32'd98; 
32'd2277: dataIn2 = 32'd74; 
32'd2278: dataIn2 = 32'd84; 
32'd2279: dataIn2 = 32'd96; 
32'd2280: dataIn2 = 32'd57; 
32'd2281: dataIn2 = 32'd43; 
32'd2282: dataIn2 = 32'd35; 
32'd2283: dataIn2 = 32'd72; 
32'd2284: dataIn2 = 32'd85; 
32'd2285: dataIn2 = 32'd63; 
32'd2286: dataIn2 = 32'd73; 
32'd2287: dataIn2 = 32'd0; 
32'd2288: dataIn2 = 32'd60; 
32'd2289: dataIn2 = 32'd30; 
32'd2290: dataIn2 = 32'd71; 
32'd2291: dataIn2 = 32'd82; 
32'd2292: dataIn2 = 32'd7; 
32'd2293: dataIn2 = 32'd70; 
32'd2294: dataIn2 = 32'd47; 
32'd2295: dataIn2 = 32'd28; 
32'd2296: dataIn2 = 32'd42; 
32'd2297: dataIn2 = 32'd52; 
32'd2298: dataIn2 = 32'd67; 
32'd2299: dataIn2 = 32'd14; 
32'd2300: dataIn2 = 32'd29; 
32'd2301: dataIn2 = 32'd56; 
32'd2302: dataIn2 = 32'd72; 
32'd2303: dataIn2 = 32'd1; 
32'd2304: dataIn2 = 32'd34; 
32'd2305: dataIn2 = 32'd85; 
32'd2306: dataIn2 = 32'd100; 
32'd2307: dataIn2 = 32'd68; 
32'd2308: dataIn2 = 32'd19; 
32'd2309: dataIn2 = 32'd27; 
32'd2310: dataIn2 = 32'd5; 
32'd2311: dataIn2 = 32'd30; 
32'd2312: dataIn2 = 32'd88; 
32'd2313: dataIn2 = 32'd50; 
32'd2314: dataIn2 = 32'd25; 
32'd2315: dataIn2 = 32'd29; 
32'd2316: dataIn2 = 32'd82; 
32'd2317: dataIn2 = 32'd15; 
32'd2318: dataIn2 = 32'd0; 
32'd2319: dataIn2 = 32'd56; 
32'd2320: dataIn2 = 32'd81; 
32'd2321: dataIn2 = 32'd87; 
32'd2322: dataIn2 = 32'd43; 
32'd2323: dataIn2 = 32'd85; 
32'd2324: dataIn2 = 32'd47; 
32'd2325: dataIn2 = 32'd54; 
32'd2326: dataIn2 = 32'd32; 
32'd2327: dataIn2 = 32'd12; 
32'd2328: dataIn2 = 32'd21; 
32'd2329: dataIn2 = 32'd58; 
32'd2330: dataIn2 = 32'd4; 
32'd2331: dataIn2 = 32'd13; 
32'd2332: dataIn2 = 32'd77; 
32'd2333: dataIn2 = 32'd21; 
32'd2334: dataIn2 = 32'd40; 
32'd2335: dataIn2 = 32'd94; 
32'd2336: dataIn2 = 32'd83; 
32'd2337: dataIn2 = 32'd39; 
32'd2338: dataIn2 = 32'd28; 
32'd2339: dataIn2 = 32'd13; 
32'd2340: dataIn2 = 32'd49; 
32'd2341: dataIn2 = 32'd72; 
32'd2342: dataIn2 = 32'd7; 
32'd2343: dataIn2 = 32'd43; 
32'd2344: dataIn2 = 32'd98; 
32'd2345: dataIn2 = 32'd98; 
32'd2346: dataIn2 = 32'd75; 
32'd2347: dataIn2 = 32'd61; 
32'd2348: dataIn2 = 32'd55; 
32'd2349: dataIn2 = 32'd13; 
32'd2350: dataIn2 = 32'd100; 
32'd2351: dataIn2 = 32'd58; 
32'd2352: dataIn2 = 32'd43; 
32'd2353: dataIn2 = 32'd23; 
32'd2354: dataIn2 = 32'd25; 
32'd2355: dataIn2 = 32'd67; 
32'd2356: dataIn2 = 32'd37; 
32'd2357: dataIn2 = 32'd30; 
32'd2358: dataIn2 = 32'd30; 
32'd2359: dataIn2 = 32'd59; 
32'd2360: dataIn2 = 32'd20; 
32'd2361: dataIn2 = 32'd55; 
32'd2362: dataIn2 = 32'd40; 
32'd2363: dataIn2 = 32'd28; 
32'd2364: dataIn2 = 32'd42; 
32'd2365: dataIn2 = 32'd46; 
32'd2366: dataIn2 = 32'd51; 
32'd2367: dataIn2 = 32'd67; 
32'd2368: dataIn2 = 32'd56; 
32'd2369: dataIn2 = 32'd51; 
32'd2370: dataIn2 = 32'd100; 
32'd2371: dataIn2 = 32'd54; 
32'd2372: dataIn2 = 32'd94; 
32'd2373: dataIn2 = 32'd65; 
32'd2374: dataIn2 = 32'd29; 
32'd2375: dataIn2 = 32'd81; 
32'd2376: dataIn2 = 32'd69; 
32'd2377: dataIn2 = 32'd6; 
32'd2378: dataIn2 = 32'd81; 
32'd2379: dataIn2 = 32'd48; 
32'd2380: dataIn2 = 32'd41; 
32'd2381: dataIn2 = 32'd20; 
32'd2382: dataIn2 = 32'd33; 
32'd2383: dataIn2 = 32'd96; 
32'd2384: dataIn2 = 32'd79; 
32'd2385: dataIn2 = 32'd54; 
32'd2386: dataIn2 = 32'd61; 
32'd2387: dataIn2 = 32'd27; 
32'd2388: dataIn2 = 32'd60; 
32'd2389: dataIn2 = 32'd80; 
32'd2390: dataIn2 = 32'd63; 
32'd2391: dataIn2 = 32'd59; 
32'd2392: dataIn2 = 32'd28; 
32'd2393: dataIn2 = 32'd84; 
32'd2394: dataIn2 = 32'd63; 
32'd2395: dataIn2 = 32'd35; 
32'd2396: dataIn2 = 32'd39; 
32'd2397: dataIn2 = 32'd44; 
32'd2398: dataIn2 = 32'd23; 
32'd2399: dataIn2 = 32'd0; 
32'd2400: dataIn2 = 32'd45; 
32'd2401: dataIn2 = 32'd78; 
32'd2402: dataIn2 = 32'd75; 
32'd2403: dataIn2 = 32'd74; 
32'd2404: dataIn2 = 32'd75; 
32'd2405: dataIn2 = 32'd6; 
32'd2406: dataIn2 = 32'd1; 
32'd2407: dataIn2 = 32'd5; 
32'd2408: dataIn2 = 32'd32; 
32'd2409: dataIn2 = 32'd20; 
32'd2410: dataIn2 = 32'd17; 
32'd2411: dataIn2 = 32'd61; 
32'd2412: dataIn2 = 32'd50; 
32'd2413: dataIn2 = 32'd8; 
32'd2414: dataIn2 = 32'd84; 
32'd2415: dataIn2 = 32'd6; 
32'd2416: dataIn2 = 32'd21; 
32'd2417: dataIn2 = 32'd70; 
32'd2418: dataIn2 = 32'd38; 
32'd2419: dataIn2 = 32'd79; 
32'd2420: dataIn2 = 32'd98; 
32'd2421: dataIn2 = 32'd26; 
32'd2422: dataIn2 = 32'd90; 
32'd2423: dataIn2 = 32'd4; 
32'd2424: dataIn2 = 32'd54; 
32'd2425: dataIn2 = 32'd42; 
32'd2426: dataIn2 = 32'd63; 
32'd2427: dataIn2 = 32'd5; 
32'd2428: dataIn2 = 32'd71; 
32'd2429: dataIn2 = 32'd20; 
32'd2430: dataIn2 = 32'd59; 
32'd2431: dataIn2 = 32'd100; 
32'd2432: dataIn2 = 32'd62; 
32'd2433: dataIn2 = 32'd100; 
32'd2434: dataIn2 = 32'd61; 
32'd2435: dataIn2 = 32'd12; 
32'd2436: dataIn2 = 32'd60; 
32'd2437: dataIn2 = 32'd75; 
32'd2438: dataIn2 = 32'd55; 
32'd2439: dataIn2 = 32'd51; 
32'd2440: dataIn2 = 32'd10; 
32'd2441: dataIn2 = 32'd9; 
32'd2442: dataIn2 = 32'd74; 
32'd2443: dataIn2 = 32'd11; 
32'd2444: dataIn2 = 32'd78; 
32'd2445: dataIn2 = 32'd21; 
32'd2446: dataIn2 = 32'd29; 
32'd2447: dataIn2 = 32'd48; 
32'd2448: dataIn2 = 32'd85; 
32'd2449: dataIn2 = 32'd53; 
32'd2450: dataIn2 = 32'd94; 
32'd2451: dataIn2 = 32'd3; 
32'd2452: dataIn2 = 32'd7; 
32'd2453: dataIn2 = 32'd44; 
32'd2454: dataIn2 = 32'd76; 
32'd2455: dataIn2 = 32'd18; 
32'd2456: dataIn2 = 32'd22; 
32'd2457: dataIn2 = 32'd93; 
32'd2458: dataIn2 = 32'd45; 
32'd2459: dataIn2 = 32'd28; 
32'd2460: dataIn2 = 32'd50; 
32'd2461: dataIn2 = 32'd44; 
32'd2462: dataIn2 = 32'd17; 
32'd2463: dataIn2 = 32'd27; 
32'd2464: dataIn2 = 32'd10; 
32'd2465: dataIn2 = 32'd61; 
32'd2466: dataIn2 = 32'd4; 
32'd2467: dataIn2 = 32'd43; 
32'd2468: dataIn2 = 32'd50; 
32'd2469: dataIn2 = 32'd39; 
32'd2470: dataIn2 = 32'd1; 
32'd2471: dataIn2 = 32'd4; 
32'd2472: dataIn2 = 32'd43; 
32'd2473: dataIn2 = 32'd34; 
32'd2474: dataIn2 = 32'd90; 
32'd2475: dataIn2 = 32'd23; 
32'd2476: dataIn2 = 32'd37; 
32'd2477: dataIn2 = 32'd43; 
32'd2478: dataIn2 = 32'd44; 
32'd2479: dataIn2 = 32'd65; 
32'd2480: dataIn2 = 32'd40; 
32'd2481: dataIn2 = 32'd69; 
32'd2482: dataIn2 = 32'd59; 
32'd2483: dataIn2 = 32'd81; 
32'd2484: dataIn2 = 32'd41; 
32'd2485: dataIn2 = 32'd14; 
32'd2486: dataIn2 = 32'd12; 
32'd2487: dataIn2 = 32'd62; 
32'd2488: dataIn2 = 32'd7; 
32'd2489: dataIn2 = 32'd86; 
32'd2490: dataIn2 = 32'd53; 
32'd2491: dataIn2 = 32'd50; 
32'd2492: dataIn2 = 32'd45; 
32'd2493: dataIn2 = 32'd38; 
32'd2494: dataIn2 = 32'd63; 
32'd2495: dataIn2 = 32'd96; 
32'd2496: dataIn2 = 32'd53; 
32'd2497: dataIn2 = 32'd65; 
32'd2498: dataIn2 = 32'd27; 
32'd2499: dataIn2 = 32'd29; 
32'd2500: dataIn2 = 32'd44; 
32'd2501: dataIn2 = 32'd1; 
32'd2502: dataIn2 = 32'd56; 
32'd2503: dataIn2 = 32'd60; 
32'd2504: dataIn2 = 32'd78; 
32'd2505: dataIn2 = 32'd90; 
32'd2506: dataIn2 = 32'd34; 
32'd2507: dataIn2 = 32'd37; 
32'd2508: dataIn2 = 32'd57; 
32'd2509: dataIn2 = 32'd55; 
32'd2510: dataIn2 = 32'd70; 
32'd2511: dataIn2 = 32'd37; 
32'd2512: dataIn2 = 32'd87; 
32'd2513: dataIn2 = 32'd28; 
32'd2514: dataIn2 = 32'd32; 
32'd2515: dataIn2 = 32'd24; 
32'd2516: dataIn2 = 32'd74; 
32'd2517: dataIn2 = 32'd58; 
32'd2518: dataIn2 = 32'd71; 
32'd2519: dataIn2 = 32'd38; 
32'd2520: dataIn2 = 32'd95; 
32'd2521: dataIn2 = 32'd4; 
32'd2522: dataIn2 = 32'd12; 
32'd2523: dataIn2 = 32'd19; 
32'd2524: dataIn2 = 32'd100; 
32'd2525: dataIn2 = 32'd84; 
32'd2526: dataIn2 = 32'd32; 
32'd2527: dataIn2 = 32'd91; 
32'd2528: dataIn2 = 32'd23; 
32'd2529: dataIn2 = 32'd93; 
32'd2530: dataIn2 = 32'd42; 
32'd2531: dataIn2 = 32'd10; 
32'd2532: dataIn2 = 32'd64; 
32'd2533: dataIn2 = 32'd31; 
32'd2534: dataIn2 = 32'd18; 
32'd2535: dataIn2 = 32'd16; 
32'd2536: dataIn2 = 32'd79; 
32'd2537: dataIn2 = 32'd73; 
32'd2538: dataIn2 = 32'd60; 
32'd2539: dataIn2 = 32'd23; 
32'd2540: dataIn2 = 32'd83; 
32'd2541: dataIn2 = 32'd5; 
32'd2542: dataIn2 = 32'd38; 
32'd2543: dataIn2 = 32'd74; 
32'd2544: dataIn2 = 32'd48; 
32'd2545: dataIn2 = 32'd99; 
32'd2546: dataIn2 = 32'd87; 
32'd2547: dataIn2 = 32'd38; 
32'd2548: dataIn2 = 32'd48; 
32'd2549: dataIn2 = 32'd96; 
32'd2550: dataIn2 = 32'd54; 
32'd2551: dataIn2 = 32'd6; 
32'd2552: dataIn2 = 32'd28; 
32'd2553: dataIn2 = 32'd15; 
32'd2554: dataIn2 = 32'd8; 
32'd2555: dataIn2 = 32'd28; 
32'd2556: dataIn2 = 32'd47; 
32'd2557: dataIn2 = 32'd100; 
32'd2558: dataIn2 = 32'd13; 
32'd2559: dataIn2 = 32'd98; 
32'd2560: dataIn2 = 32'd83; 
32'd2561: dataIn2 = 32'd6; 
32'd2562: dataIn2 = 32'd10; 
32'd2563: dataIn2 = 32'd29; 
32'd2564: dataIn2 = 32'd100; 
32'd2565: dataIn2 = 32'd80; 
32'd2566: dataIn2 = 32'd80; 
32'd2567: dataIn2 = 32'd76; 
32'd2568: dataIn2 = 32'd38; 
32'd2569: dataIn2 = 32'd94; 
32'd2570: dataIn2 = 32'd95; 
32'd2571: dataIn2 = 32'd90; 
32'd2572: dataIn2 = 32'd21; 
32'd2573: dataIn2 = 32'd99; 
32'd2574: dataIn2 = 32'd21; 
32'd2575: dataIn2 = 32'd92; 
32'd2576: dataIn2 = 32'd25; 
32'd2577: dataIn2 = 32'd33; 
32'd2578: dataIn2 = 32'd72; 
32'd2579: dataIn2 = 32'd53; 
32'd2580: dataIn2 = 32'd23; 
32'd2581: dataIn2 = 32'd67; 
32'd2582: dataIn2 = 32'd43; 
32'd2583: dataIn2 = 32'd21; 
32'd2584: dataIn2 = 32'd6; 
32'd2585: dataIn2 = 32'd71; 
32'd2586: dataIn2 = 32'd68; 
32'd2587: dataIn2 = 32'd60; 
32'd2588: dataIn2 = 32'd77; 
32'd2589: dataIn2 = 32'd82; 
32'd2590: dataIn2 = 32'd27; 
32'd2591: dataIn2 = 32'd32; 
32'd2592: dataIn2 = 32'd95; 
32'd2593: dataIn2 = 32'd99; 
32'd2594: dataIn2 = 32'd77; 
32'd2595: dataIn2 = 32'd46; 
32'd2596: dataIn2 = 32'd94; 
32'd2597: dataIn2 = 32'd34; 
32'd2598: dataIn2 = 32'd20; 
32'd2599: dataIn2 = 32'd7; 
32'd2600: dataIn2 = 32'd12; 
32'd2601: dataIn2 = 32'd99; 
32'd2602: dataIn2 = 32'd62; 
32'd2603: dataIn2 = 32'd47; 
32'd2604: dataIn2 = 32'd64; 
32'd2605: dataIn2 = 32'd20; 
32'd2606: dataIn2 = 32'd96; 
32'd2607: dataIn2 = 32'd13; 
32'd2608: dataIn2 = 32'd75; 
32'd2609: dataIn2 = 32'd32; 
32'd2610: dataIn2 = 32'd84; 
32'd2611: dataIn2 = 32'd57; 
32'd2612: dataIn2 = 32'd2; 
32'd2613: dataIn2 = 32'd67; 
32'd2614: dataIn2 = 32'd10; 
32'd2615: dataIn2 = 32'd53; 
32'd2616: dataIn2 = 32'd99; 
32'd2617: dataIn2 = 32'd8; 
32'd2618: dataIn2 = 32'd38; 
32'd2619: dataIn2 = 32'd62; 
32'd2620: dataIn2 = 32'd95; 
32'd2621: dataIn2 = 32'd82; 
32'd2622: dataIn2 = 32'd86; 
32'd2623: dataIn2 = 32'd45; 
32'd2624: dataIn2 = 32'd95; 
32'd2625: dataIn2 = 32'd22; 
32'd2626: dataIn2 = 32'd46; 
32'd2627: dataIn2 = 32'd35; 
32'd2628: dataIn2 = 32'd42; 
32'd2629: dataIn2 = 32'd62; 
32'd2630: dataIn2 = 32'd93; 
32'd2631: dataIn2 = 32'd34; 
32'd2632: dataIn2 = 32'd19; 
32'd2633: dataIn2 = 32'd11; 
32'd2634: dataIn2 = 32'd29; 
32'd2635: dataIn2 = 32'd83; 
32'd2636: dataIn2 = 32'd21; 
32'd2637: dataIn2 = 32'd96; 
32'd2638: dataIn2 = 32'd30; 
32'd2639: dataIn2 = 32'd17; 
32'd2640: dataIn2 = 32'd17; 
32'd2641: dataIn2 = 32'd39; 
32'd2642: dataIn2 = 32'd1; 
32'd2643: dataIn2 = 32'd83; 
32'd2644: dataIn2 = 32'd79; 
32'd2645: dataIn2 = 32'd72; 
32'd2646: dataIn2 = 32'd56; 
32'd2647: dataIn2 = 32'd72; 
32'd2648: dataIn2 = 32'd93; 
32'd2649: dataIn2 = 32'd44; 
32'd2650: dataIn2 = 32'd69; 
32'd2651: dataIn2 = 32'd72; 
32'd2652: dataIn2 = 32'd62; 
32'd2653: dataIn2 = 32'd53; 
32'd2654: dataIn2 = 32'd41; 
32'd2655: dataIn2 = 32'd18; 
32'd2656: dataIn2 = 32'd19; 
32'd2657: dataIn2 = 32'd100; 
32'd2658: dataIn2 = 32'd74; 
32'd2659: dataIn2 = 32'd70; 
32'd2660: dataIn2 = 32'd27; 
32'd2661: dataIn2 = 32'd30; 
32'd2662: dataIn2 = 32'd30; 
32'd2663: dataIn2 = 32'd57; 
32'd2664: dataIn2 = 32'd15; 
32'd2665: dataIn2 = 32'd76; 
32'd2666: dataIn2 = 32'd46; 
32'd2667: dataIn2 = 32'd84; 
32'd2668: dataIn2 = 32'd76; 
32'd2669: dataIn2 = 32'd7; 
32'd2670: dataIn2 = 32'd41; 
32'd2671: dataIn2 = 32'd82; 
32'd2672: dataIn2 = 32'd11; 
32'd2673: dataIn2 = 32'd50; 
32'd2674: dataIn2 = 32'd33; 
32'd2675: dataIn2 = 32'd28; 
32'd2676: dataIn2 = 32'd55; 
32'd2677: dataIn2 = 32'd57; 
32'd2678: dataIn2 = 32'd65; 
32'd2679: dataIn2 = 32'd77; 
32'd2680: dataIn2 = 32'd0; 
32'd2681: dataIn2 = 32'd39; 
32'd2682: dataIn2 = 32'd57; 
32'd2683: dataIn2 = 32'd50; 
32'd2684: dataIn2 = 32'd27; 
32'd2685: dataIn2 = 32'd3; 
32'd2686: dataIn2 = 32'd62; 
32'd2687: dataIn2 = 32'd29; 
32'd2688: dataIn2 = 32'd91; 
32'd2689: dataIn2 = 32'd68; 
32'd2690: dataIn2 = 32'd97; 
32'd2691: dataIn2 = 32'd86; 
32'd2692: dataIn2 = 32'd54; 
32'd2693: dataIn2 = 32'd42; 
32'd2694: dataIn2 = 32'd60; 
32'd2695: dataIn2 = 32'd32; 
32'd2696: dataIn2 = 32'd100; 
32'd2697: dataIn2 = 32'd69; 
32'd2698: dataIn2 = 32'd58; 
32'd2699: dataIn2 = 32'd69; 
32'd2700: dataIn2 = 32'd76; 
32'd2701: dataIn2 = 32'd14; 
32'd2702: dataIn2 = 32'd81; 
32'd2703: dataIn2 = 32'd39; 
32'd2704: dataIn2 = 32'd44; 
32'd2705: dataIn2 = 32'd47; 
32'd2706: dataIn2 = 32'd77; 
32'd2707: dataIn2 = 32'd17; 
32'd2708: dataIn2 = 32'd60; 
32'd2709: dataIn2 = 32'd45; 
32'd2710: dataIn2 = 32'd5; 
32'd2711: dataIn2 = 32'd40; 
32'd2712: dataIn2 = 32'd75; 
32'd2713: dataIn2 = 32'd18; 
32'd2714: dataIn2 = 32'd23; 
32'd2715: dataIn2 = 32'd19; 
32'd2716: dataIn2 = 32'd52; 
32'd2717: dataIn2 = 32'd80; 
32'd2718: dataIn2 = 32'd93; 
32'd2719: dataIn2 = 32'd12; 
32'd2720: dataIn2 = 32'd85; 
32'd2721: dataIn2 = 32'd59; 
32'd2722: dataIn2 = 32'd32; 
32'd2723: dataIn2 = 32'd12; 
32'd2724: dataIn2 = 32'd99; 
32'd2725: dataIn2 = 32'd58; 
32'd2726: dataIn2 = 32'd30; 
32'd2727: dataIn2 = 32'd56; 
32'd2728: dataIn2 = 32'd27; 
32'd2729: dataIn2 = 32'd50; 
32'd2730: dataIn2 = 32'd12; 
32'd2731: dataIn2 = 32'd70; 
32'd2732: dataIn2 = 32'd88; 
32'd2733: dataIn2 = 32'd13; 
32'd2734: dataIn2 = 32'd23; 
32'd2735: dataIn2 = 32'd46; 
32'd2736: dataIn2 = 32'd43; 
32'd2737: dataIn2 = 32'd83; 
32'd2738: dataIn2 = 32'd97; 
32'd2739: dataIn2 = 32'd62; 
32'd2740: dataIn2 = 32'd70; 
32'd2741: dataIn2 = 32'd85; 
32'd2742: dataIn2 = 32'd13; 
32'd2743: dataIn2 = 32'd43; 
32'd2744: dataIn2 = 32'd10; 
32'd2745: dataIn2 = 32'd19; 
32'd2746: dataIn2 = 32'd4; 
32'd2747: dataIn2 = 32'd82; 
32'd2748: dataIn2 = 32'd35; 
32'd2749: dataIn2 = 32'd80; 
32'd2750: dataIn2 = 32'd40; 
32'd2751: dataIn2 = 32'd58; 
32'd2752: dataIn2 = 32'd42; 
32'd2753: dataIn2 = 32'd72; 
32'd2754: dataIn2 = 32'd38; 
32'd2755: dataIn2 = 32'd49; 
32'd2756: dataIn2 = 32'd43; 
32'd2757: dataIn2 = 32'd29; 
32'd2758: dataIn2 = 32'd59; 
32'd2759: dataIn2 = 32'd26; 
32'd2760: dataIn2 = 32'd57; 
32'd2761: dataIn2 = 32'd81; 
32'd2762: dataIn2 = 32'd89; 
32'd2763: dataIn2 = 32'd19; 
32'd2764: dataIn2 = 32'd50; 
32'd2765: dataIn2 = 32'd69; 
32'd2766: dataIn2 = 32'd74; 
32'd2767: dataIn2 = 32'd99; 
32'd2768: dataIn2 = 32'd68; 
32'd2769: dataIn2 = 32'd2; 
32'd2770: dataIn2 = 32'd78; 
32'd2771: dataIn2 = 32'd91; 
32'd2772: dataIn2 = 32'd70; 
32'd2773: dataIn2 = 32'd72; 
32'd2774: dataIn2 = 32'd57; 
32'd2775: dataIn2 = 32'd42; 
32'd2776: dataIn2 = 32'd96; 
32'd2777: dataIn2 = 32'd62; 
32'd2778: dataIn2 = 32'd11; 
32'd2779: dataIn2 = 32'd88; 
32'd2780: dataIn2 = 32'd33; 
32'd2781: dataIn2 = 32'd82; 
32'd2782: dataIn2 = 32'd11; 
32'd2783: dataIn2 = 32'd22; 
32'd2784: dataIn2 = 32'd20; 
32'd2785: dataIn2 = 32'd35; 
32'd2786: dataIn2 = 32'd4; 
32'd2787: dataIn2 = 32'd25; 
32'd2788: dataIn2 = 32'd2; 
32'd2789: dataIn2 = 32'd82; 
32'd2790: dataIn2 = 32'd42; 
32'd2791: dataIn2 = 32'd48; 
32'd2792: dataIn2 = 32'd89; 
32'd2793: dataIn2 = 32'd49; 
32'd2794: dataIn2 = 32'd39; 
32'd2795: dataIn2 = 32'd30; 
32'd2796: dataIn2 = 32'd37; 
32'd2797: dataIn2 = 32'd73; 
32'd2798: dataIn2 = 32'd13; 
32'd2799: dataIn2 = 32'd16; 
32'd2800: dataIn2 = 32'd73; 
32'd2801: dataIn2 = 32'd51; 
32'd2802: dataIn2 = 32'd93; 
32'd2803: dataIn2 = 32'd52; 
32'd2804: dataIn2 = 32'd43; 
32'd2805: dataIn2 = 32'd36; 
32'd2806: dataIn2 = 32'd9; 
32'd2807: dataIn2 = 32'd20; 
32'd2808: dataIn2 = 32'd66; 
32'd2809: dataIn2 = 32'd21; 
32'd2810: dataIn2 = 32'd59; 
32'd2811: dataIn2 = 32'd51; 
32'd2812: dataIn2 = 32'd34; 
32'd2813: dataIn2 = 32'd15; 
32'd2814: dataIn2 = 32'd97; 
32'd2815: dataIn2 = 32'd48; 
32'd2816: dataIn2 = 32'd14; 
32'd2817: dataIn2 = 32'd18; 
32'd2818: dataIn2 = 32'd64; 
32'd2819: dataIn2 = 32'd84; 
32'd2820: dataIn2 = 32'd14; 
32'd2821: dataIn2 = 32'd17; 
32'd2822: dataIn2 = 32'd47; 
32'd2823: dataIn2 = 32'd28; 
32'd2824: dataIn2 = 32'd29; 
32'd2825: dataIn2 = 32'd97; 
32'd2826: dataIn2 = 32'd37; 
32'd2827: dataIn2 = 32'd65; 
32'd2828: dataIn2 = 32'd42; 
32'd2829: dataIn2 = 32'd87; 
32'd2830: dataIn2 = 32'd50; 
32'd2831: dataIn2 = 32'd81; 
32'd2832: dataIn2 = 32'd80; 
32'd2833: dataIn2 = 32'd65; 
32'd2834: dataIn2 = 32'd49; 
32'd2835: dataIn2 = 32'd47; 
32'd2836: dataIn2 = 32'd87; 
32'd2837: dataIn2 = 32'd96; 
32'd2838: dataIn2 = 32'd11; 
32'd2839: dataIn2 = 32'd70; 
32'd2840: dataIn2 = 32'd71; 
32'd2841: dataIn2 = 32'd55; 
32'd2842: dataIn2 = 32'd17; 
32'd2843: dataIn2 = 32'd47; 
32'd2844: dataIn2 = 32'd35; 
32'd2845: dataIn2 = 32'd76; 
32'd2846: dataIn2 = 32'd83; 
32'd2847: dataIn2 = 32'd19; 
32'd2848: dataIn2 = 32'd84; 
32'd2849: dataIn2 = 32'd48; 
32'd2850: dataIn2 = 32'd94; 
32'd2851: dataIn2 = 32'd6; 
32'd2852: dataIn2 = 32'd27; 
32'd2853: dataIn2 = 32'd53; 
32'd2854: dataIn2 = 32'd76; 
32'd2855: dataIn2 = 32'd75; 
32'd2856: dataIn2 = 32'd53; 
32'd2857: dataIn2 = 32'd64; 
32'd2858: dataIn2 = 32'd32; 
32'd2859: dataIn2 = 32'd29; 
32'd2860: dataIn2 = 32'd49; 
32'd2861: dataIn2 = 32'd74; 
32'd2862: dataIn2 = 32'd66; 
32'd2863: dataIn2 = 32'd56; 
32'd2864: dataIn2 = 32'd74; 
32'd2865: dataIn2 = 32'd4; 
32'd2866: dataIn2 = 32'd93; 
32'd2867: dataIn2 = 32'd48; 
32'd2868: dataIn2 = 32'd1; 
32'd2869: dataIn2 = 32'd13; 
32'd2870: dataIn2 = 32'd78; 
32'd2871: dataIn2 = 32'd22; 
32'd2872: dataIn2 = 32'd86; 
32'd2873: dataIn2 = 32'd50; 
32'd2874: dataIn2 = 32'd49; 
32'd2875: dataIn2 = 32'd36; 
32'd2876: dataIn2 = 32'd22; 
32'd2877: dataIn2 = 32'd36; 
32'd2878: dataIn2 = 32'd94; 
32'd2879: dataIn2 = 32'd32; 
32'd2880: dataIn2 = 32'd21; 
32'd2881: dataIn2 = 32'd42; 
32'd2882: dataIn2 = 32'd5; 
32'd2883: dataIn2 = 32'd67; 
32'd2884: dataIn2 = 32'd92; 
32'd2885: dataIn2 = 32'd63; 
32'd2886: dataIn2 = 32'd71; 
32'd2887: dataIn2 = 32'd42; 
32'd2888: dataIn2 = 32'd84; 
32'd2889: dataIn2 = 32'd16; 
32'd2890: dataIn2 = 32'd41; 
32'd2891: dataIn2 = 32'd56; 
32'd2892: dataIn2 = 32'd97; 
32'd2893: dataIn2 = 32'd44; 
32'd2894: dataIn2 = 32'd32; 
32'd2895: dataIn2 = 32'd51; 
32'd2896: dataIn2 = 32'd66; 
32'd2897: dataIn2 = 32'd33; 
32'd2898: dataIn2 = 32'd19; 
32'd2899: dataIn2 = 32'd73; 
32'd2900: dataIn2 = 32'd65; 
32'd2901: dataIn2 = 32'd97; 
32'd2902: dataIn2 = 32'd25; 
32'd2903: dataIn2 = 32'd8; 
32'd2904: dataIn2 = 32'd95; 
32'd2905: dataIn2 = 32'd13; 
32'd2906: dataIn2 = 32'd17; 
32'd2907: dataIn2 = 32'd50; 
32'd2908: dataIn2 = 32'd23; 
32'd2909: dataIn2 = 32'd59; 
32'd2910: dataIn2 = 32'd69; 
32'd2911: dataIn2 = 32'd62; 
32'd2912: dataIn2 = 32'd31; 
32'd2913: dataIn2 = 32'd46; 
32'd2914: dataIn2 = 32'd33; 
32'd2915: dataIn2 = 32'd49; 
32'd2916: dataIn2 = 32'd10; 
32'd2917: dataIn2 = 32'd64; 
32'd2918: dataIn2 = 32'd85; 
32'd2919: dataIn2 = 32'd39; 
32'd2920: dataIn2 = 32'd15; 
32'd2921: dataIn2 = 32'd36; 
32'd2922: dataIn2 = 32'd63; 
32'd2923: dataIn2 = 32'd24; 
32'd2924: dataIn2 = 32'd95; 
32'd2925: dataIn2 = 32'd35; 
32'd2926: dataIn2 = 32'd34; 
32'd2927: dataIn2 = 32'd59; 
32'd2928: dataIn2 = 32'd53; 
32'd2929: dataIn2 = 32'd44; 
32'd2930: dataIn2 = 32'd55; 
32'd2931: dataIn2 = 32'd71; 
32'd2932: dataIn2 = 32'd70; 
32'd2933: dataIn2 = 32'd99; 
32'd2934: dataIn2 = 32'd42; 
32'd2935: dataIn2 = 32'd32; 
32'd2936: dataIn2 = 32'd67; 
32'd2937: dataIn2 = 32'd56; 
32'd2938: dataIn2 = 32'd83; 
32'd2939: dataIn2 = 32'd53; 
32'd2940: dataIn2 = 32'd95; 
32'd2941: dataIn2 = 32'd38; 
32'd2942: dataIn2 = 32'd33; 
32'd2943: dataIn2 = 32'd54; 
32'd2944: dataIn2 = 32'd19; 
32'd2945: dataIn2 = 32'd8; 
32'd2946: dataIn2 = 32'd49; 
32'd2947: dataIn2 = 32'd52; 
32'd2948: dataIn2 = 32'd58; 
32'd2949: dataIn2 = 32'd64; 
32'd2950: dataIn2 = 32'd34; 
32'd2951: dataIn2 = 32'd5; 
32'd2952: dataIn2 = 32'd94; 
32'd2953: dataIn2 = 32'd76; 
32'd2954: dataIn2 = 32'd15; 
32'd2955: dataIn2 = 32'd97; 
32'd2956: dataIn2 = 32'd49; 
32'd2957: dataIn2 = 32'd90; 
32'd2958: dataIn2 = 32'd68; 
32'd2959: dataIn2 = 32'd36; 
32'd2960: dataIn2 = 32'd94; 
32'd2961: dataIn2 = 32'd50; 
32'd2962: dataIn2 = 32'd65; 
32'd2963: dataIn2 = 32'd35; 
32'd2964: dataIn2 = 32'd7; 
32'd2965: dataIn2 = 32'd68; 
32'd2966: dataIn2 = 32'd75; 
32'd2967: dataIn2 = 32'd41; 
32'd2968: dataIn2 = 32'd52; 
32'd2969: dataIn2 = 32'd38; 
32'd2970: dataIn2 = 32'd16; 
32'd2971: dataIn2 = 32'd100; 
32'd2972: dataIn2 = 32'd72; 
32'd2973: dataIn2 = 32'd68; 
32'd2974: dataIn2 = 32'd20; 
32'd2975: dataIn2 = 32'd6; 
32'd2976: dataIn2 = 32'd96; 
32'd2977: dataIn2 = 32'd31; 
32'd2978: dataIn2 = 32'd92; 
32'd2979: dataIn2 = 32'd77; 
32'd2980: dataIn2 = 32'd16; 
32'd2981: dataIn2 = 32'd23; 
32'd2982: dataIn2 = 32'd92; 
32'd2983: dataIn2 = 32'd83; 
32'd2984: dataIn2 = 32'd93; 
32'd2985: dataIn2 = 32'd38; 
32'd2986: dataIn2 = 32'd27; 
32'd2987: dataIn2 = 32'd98; 
32'd2988: dataIn2 = 32'd2; 
32'd2989: dataIn2 = 32'd46; 
32'd2990: dataIn2 = 32'd50; 
32'd2991: dataIn2 = 32'd1; 
32'd2992: dataIn2 = 32'd82; 
32'd2993: dataIn2 = 32'd39; 
32'd2994: dataIn2 = 32'd50; 
32'd2995: dataIn2 = 32'd13; 
32'd2996: dataIn2 = 32'd16; 
32'd2997: dataIn2 = 32'd71; 
32'd2998: dataIn2 = 32'd11; 
32'd2999: dataIn2 = 32'd22; 
32'd3000: dataIn2 = 32'd20; 
32'd3001: dataIn2 = 32'd68; 
32'd3002: dataIn2 = 32'd84; 
32'd3003: dataIn2 = 32'd56; 
32'd3004: dataIn2 = 32'd71; 
32'd3005: dataIn2 = 32'd95; 
32'd3006: dataIn2 = 32'd28; 
32'd3007: dataIn2 = 32'd19; 
32'd3008: dataIn2 = 32'd7; 
32'd3009: dataIn2 = 32'd26; 
32'd3010: dataIn2 = 32'd49; 
32'd3011: dataIn2 = 32'd12; 
32'd3012: dataIn2 = 32'd32; 
32'd3013: dataIn2 = 32'd50; 
32'd3014: dataIn2 = 32'd22; 
32'd3015: dataIn2 = 32'd95; 
32'd3016: dataIn2 = 32'd63; 
32'd3017: dataIn2 = 32'd42; 
32'd3018: dataIn2 = 32'd6; 
32'd3019: dataIn2 = 32'd14; 
32'd3020: dataIn2 = 32'd98; 
32'd3021: dataIn2 = 32'd11; 
32'd3022: dataIn2 = 32'd1; 
32'd3023: dataIn2 = 32'd41; 
32'd3024: dataIn2 = 32'd28; 
32'd3025: dataIn2 = 32'd76; 
32'd3026: dataIn2 = 32'd56; 
32'd3027: dataIn2 = 32'd86; 
32'd3028: dataIn2 = 32'd79; 
32'd3029: dataIn2 = 32'd91; 
32'd3030: dataIn2 = 32'd0; 
32'd3031: dataIn2 = 32'd40; 
32'd3032: dataIn2 = 32'd43; 
32'd3033: dataIn2 = 32'd45; 
32'd3034: dataIn2 = 32'd67; 
32'd3035: dataIn2 = 32'd30; 
32'd3036: dataIn2 = 32'd72; 
32'd3037: dataIn2 = 32'd27; 
32'd3038: dataIn2 = 32'd15; 
32'd3039: dataIn2 = 32'd52; 
32'd3040: dataIn2 = 32'd56; 
32'd3041: dataIn2 = 32'd18; 
32'd3042: dataIn2 = 32'd74; 
32'd3043: dataIn2 = 32'd76; 
32'd3044: dataIn2 = 32'd28; 
32'd3045: dataIn2 = 32'd80; 
32'd3046: dataIn2 = 32'd79; 
32'd3047: dataIn2 = 32'd51; 
32'd3048: dataIn2 = 32'd17; 
32'd3049: dataIn2 = 32'd81; 
32'd3050: dataIn2 = 32'd56; 
32'd3051: dataIn2 = 32'd55; 
32'd3052: dataIn2 = 32'd4; 
32'd3053: dataIn2 = 32'd34; 
32'd3054: dataIn2 = 32'd34; 
32'd3055: dataIn2 = 32'd43; 
32'd3056: dataIn2 = 32'd74; 
32'd3057: dataIn2 = 32'd100; 
32'd3058: dataIn2 = 32'd35; 
32'd3059: dataIn2 = 32'd23; 
32'd3060: dataIn2 = 32'd33; 
32'd3061: dataIn2 = 32'd39; 
32'd3062: dataIn2 = 32'd26; 
32'd3063: dataIn2 = 32'd53; 
32'd3064: dataIn2 = 32'd52; 
32'd3065: dataIn2 = 32'd57; 
32'd3066: dataIn2 = 32'd47; 
32'd3067: dataIn2 = 32'd38; 
32'd3068: dataIn2 = 32'd56; 
32'd3069: dataIn2 = 32'd4; 
32'd3070: dataIn2 = 32'd19; 
32'd3071: dataIn2 = 32'd51; 
32'd3072: dataIn2 = 32'd21; 
32'd3073: dataIn2 = 32'd44; 
32'd3074: dataIn2 = 32'd49; 
32'd3075: dataIn2 = 32'd88; 
32'd3076: dataIn2 = 32'd76; 
32'd3077: dataIn2 = 32'd61; 
32'd3078: dataIn2 = 32'd32; 
32'd3079: dataIn2 = 32'd60; 
32'd3080: dataIn2 = 32'd83; 
32'd3081: dataIn2 = 32'd75; 
32'd3082: dataIn2 = 32'd100; 
32'd3083: dataIn2 = 32'd64; 
32'd3084: dataIn2 = 32'd36; 
32'd3085: dataIn2 = 32'd2; 
32'd3086: dataIn2 = 32'd39; 
32'd3087: dataIn2 = 32'd17; 
32'd3088: dataIn2 = 32'd98; 
32'd3089: dataIn2 = 32'd79; 
32'd3090: dataIn2 = 32'd4; 
32'd3091: dataIn2 = 32'd0; 
32'd3092: dataIn2 = 32'd57; 
32'd3093: dataIn2 = 32'd19; 
32'd3094: dataIn2 = 32'd20; 
32'd3095: dataIn2 = 32'd30; 
32'd3096: dataIn2 = 32'd53; 
32'd3097: dataIn2 = 32'd70; 
32'd3098: dataIn2 = 32'd36; 
32'd3099: dataIn2 = 32'd33; 
32'd3100: dataIn2 = 32'd57; 
32'd3101: dataIn2 = 32'd90; 
32'd3102: dataIn2 = 32'd42; 
32'd3103: dataIn2 = 32'd81; 
32'd3104: dataIn2 = 32'd42; 
32'd3105: dataIn2 = 32'd26; 
32'd3106: dataIn2 = 32'd50; 
32'd3107: dataIn2 = 32'd72; 
32'd3108: dataIn2 = 32'd75; 
32'd3109: dataIn2 = 32'd22; 
32'd3110: dataIn2 = 32'd23; 
32'd3111: dataIn2 = 32'd29; 
32'd3112: dataIn2 = 32'd58; 
32'd3113: dataIn2 = 32'd45; 
32'd3114: dataIn2 = 32'd45; 
32'd3115: dataIn2 = 32'd30; 
32'd3116: dataIn2 = 32'd56; 
32'd3117: dataIn2 = 32'd19; 
32'd3118: dataIn2 = 32'd92; 
32'd3119: dataIn2 = 32'd45; 
32'd3120: dataIn2 = 32'd80; 
32'd3121: dataIn2 = 32'd60; 
32'd3122: dataIn2 = 32'd89; 
32'd3123: dataIn2 = 32'd79; 
32'd3124: dataIn2 = 32'd20; 
32'd3125: dataIn2 = 32'd100; 
32'd3126: dataIn2 = 32'd45; 
32'd3127: dataIn2 = 32'd95; 
32'd3128: dataIn2 = 32'd36; 
32'd3129: dataIn2 = 32'd53; 
32'd3130: dataIn2 = 32'd35; 
32'd3131: dataIn2 = 32'd85; 
32'd3132: dataIn2 = 32'd81; 
32'd3133: dataIn2 = 32'd51; 
32'd3134: dataIn2 = 32'd17; 
32'd3135: dataIn2 = 32'd100; 
32'd3136: dataIn2 = 32'd29; 
32'd3137: dataIn2 = 32'd20; 
32'd3138: dataIn2 = 32'd47; 
32'd3139: dataIn2 = 32'd46; 
32'd3140: dataIn2 = 32'd82; 
32'd3141: dataIn2 = 32'd32; 
32'd3142: dataIn2 = 32'd61; 
32'd3143: dataIn2 = 32'd25; 
32'd3144: dataIn2 = 32'd94; 
32'd3145: dataIn2 = 32'd32; 
32'd3146: dataIn2 = 32'd98; 
32'd3147: dataIn2 = 32'd21; 
32'd3148: dataIn2 = 32'd93; 
32'd3149: dataIn2 = 32'd95; 
32'd3150: dataIn2 = 32'd70; 
32'd3151: dataIn2 = 32'd37; 
32'd3152: dataIn2 = 32'd92; 
32'd3153: dataIn2 = 32'd6; 
32'd3154: dataIn2 = 32'd56; 
32'd3155: dataIn2 = 32'd37; 
32'd3156: dataIn2 = 32'd54; 
32'd3157: dataIn2 = 32'd19; 
32'd3158: dataIn2 = 32'd19; 
32'd3159: dataIn2 = 32'd12; 
32'd3160: dataIn2 = 32'd44; 
32'd3161: dataIn2 = 32'd0; 
32'd3162: dataIn2 = 32'd36; 
32'd3163: dataIn2 = 32'd70; 
32'd3164: dataIn2 = 32'd17; 
32'd3165: dataIn2 = 32'd5; 
32'd3166: dataIn2 = 32'd32; 
32'd3167: dataIn2 = 32'd80; 
32'd3168: dataIn2 = 32'd17; 
32'd3169: dataIn2 = 32'd58; 
32'd3170: dataIn2 = 32'd41; 
32'd3171: dataIn2 = 32'd76; 
32'd3172: dataIn2 = 32'd49; 
32'd3173: dataIn2 = 32'd6; 
32'd3174: dataIn2 = 32'd97; 
32'd3175: dataIn2 = 32'd84; 
32'd3176: dataIn2 = 32'd31; 
32'd3177: dataIn2 = 32'd58; 
32'd3178: dataIn2 = 32'd81; 
32'd3179: dataIn2 = 32'd58; 
32'd3180: dataIn2 = 32'd97; 
32'd3181: dataIn2 = 32'd64; 
32'd3182: dataIn2 = 32'd13; 
32'd3183: dataIn2 = 32'd80; 
32'd3184: dataIn2 = 32'd88; 
32'd3185: dataIn2 = 32'd18; 
32'd3186: dataIn2 = 32'd56; 
32'd3187: dataIn2 = 32'd96; 
32'd3188: dataIn2 = 32'd52; 
32'd3189: dataIn2 = 32'd71; 
32'd3190: dataIn2 = 32'd25; 
32'd3191: dataIn2 = 32'd51; 
32'd3192: dataIn2 = 32'd15; 
32'd3193: dataIn2 = 32'd7; 
32'd3194: dataIn2 = 32'd95; 
32'd3195: dataIn2 = 32'd4; 
32'd3196: dataIn2 = 32'd88; 
32'd3197: dataIn2 = 32'd62; 
32'd3198: dataIn2 = 32'd7; 
32'd3199: dataIn2 = 32'd18; 
32'd3200: dataIn2 = 32'd62; 
32'd3201: dataIn2 = 32'd93; 
32'd3202: dataIn2 = 32'd13; 
32'd3203: dataIn2 = 32'd51; 
32'd3204: dataIn2 = 32'd85; 
32'd3205: dataIn2 = 32'd6; 
32'd3206: dataIn2 = 32'd91; 
32'd3207: dataIn2 = 32'd30; 
32'd3208: dataIn2 = 32'd18; 
32'd3209: dataIn2 = 32'd12; 
32'd3210: dataIn2 = 32'd94; 
32'd3211: dataIn2 = 32'd50; 
32'd3212: dataIn2 = 32'd31; 
32'd3213: dataIn2 = 32'd5; 
32'd3214: dataIn2 = 32'd2; 
32'd3215: dataIn2 = 32'd67; 
32'd3216: dataIn2 = 32'd76; 
32'd3217: dataIn2 = 32'd11; 
32'd3218: dataIn2 = 32'd13; 
32'd3219: dataIn2 = 32'd3; 
32'd3220: dataIn2 = 32'd76; 
32'd3221: dataIn2 = 32'd91; 
32'd3222: dataIn2 = 32'd82; 
32'd3223: dataIn2 = 32'd4; 
32'd3224: dataIn2 = 32'd51; 
32'd3225: dataIn2 = 32'd50; 
32'd3226: dataIn2 = 32'd58; 
32'd3227: dataIn2 = 32'd91; 
32'd3228: dataIn2 = 32'd49; 
32'd3229: dataIn2 = 32'd60; 
32'd3230: dataIn2 = 32'd51; 
32'd3231: dataIn2 = 32'd5; 
32'd3232: dataIn2 = 32'd77; 
32'd3233: dataIn2 = 32'd60; 
32'd3234: dataIn2 = 32'd13; 
32'd3235: dataIn2 = 32'd37; 
32'd3236: dataIn2 = 32'd72; 
32'd3237: dataIn2 = 32'd48; 
32'd3238: dataIn2 = 32'd86; 
32'd3239: dataIn2 = 32'd4; 
32'd3240: dataIn2 = 32'd36; 
32'd3241: dataIn2 = 32'd86; 
32'd3242: dataIn2 = 32'd15; 
32'd3243: dataIn2 = 32'd51; 
32'd3244: dataIn2 = 32'd5; 
32'd3245: dataIn2 = 32'd32; 
32'd3246: dataIn2 = 32'd98; 
32'd3247: dataIn2 = 32'd59; 
32'd3248: dataIn2 = 32'd5; 
32'd3249: dataIn2 = 32'd23; 
32'd3250: dataIn2 = 32'd81; 
32'd3251: dataIn2 = 32'd73; 
32'd3252: dataIn2 = 32'd82; 
32'd3253: dataIn2 = 32'd68; 
32'd3254: dataIn2 = 32'd29; 
32'd3255: dataIn2 = 32'd0; 
32'd3256: dataIn2 = 32'd12; 
32'd3257: dataIn2 = 32'd81; 
32'd3258: dataIn2 = 32'd17; 
32'd3259: dataIn2 = 32'd24; 
32'd3260: dataIn2 = 32'd82; 
32'd3261: dataIn2 = 32'd29; 
32'd3262: dataIn2 = 32'd3; 
32'd3263: dataIn2 = 32'd97; 
32'd3264: dataIn2 = 32'd63; 
32'd3265: dataIn2 = 32'd73; 
32'd3266: dataIn2 = 32'd17; 
32'd3267: dataIn2 = 32'd86; 
32'd3268: dataIn2 = 32'd53; 
32'd3269: dataIn2 = 32'd66; 
32'd3270: dataIn2 = 32'd62; 
32'd3271: dataIn2 = 32'd2; 
32'd3272: dataIn2 = 32'd63; 
32'd3273: dataIn2 = 32'd67; 
32'd3274: dataIn2 = 32'd27; 
32'd3275: dataIn2 = 32'd7; 
32'd3276: dataIn2 = 32'd53; 
32'd3277: dataIn2 = 32'd85; 
32'd3278: dataIn2 = 32'd64; 
32'd3279: dataIn2 = 32'd62; 
32'd3280: dataIn2 = 32'd93; 
32'd3281: dataIn2 = 32'd0; 
32'd3282: dataIn2 = 32'd58; 
32'd3283: dataIn2 = 32'd78; 
32'd3284: dataIn2 = 32'd0; 
32'd3285: dataIn2 = 32'd16; 
32'd3286: dataIn2 = 32'd32; 
32'd3287: dataIn2 = 32'd95; 
32'd3288: dataIn2 = 32'd79; 
32'd3289: dataIn2 = 32'd63; 
32'd3290: dataIn2 = 32'd38; 
32'd3291: dataIn2 = 32'd31; 
32'd3292: dataIn2 = 32'd59; 
32'd3293: dataIn2 = 32'd64; 
32'd3294: dataIn2 = 32'd16; 
32'd3295: dataIn2 = 32'd95; 
32'd3296: dataIn2 = 32'd19; 
32'd3297: dataIn2 = 32'd42; 
32'd3298: dataIn2 = 32'd93; 
32'd3299: dataIn2 = 32'd68; 
32'd3300: dataIn2 = 32'd36; 
32'd3301: dataIn2 = 32'd36; 
32'd3302: dataIn2 = 32'd75; 
32'd3303: dataIn2 = 32'd89; 
32'd3304: dataIn2 = 32'd47; 
32'd3305: dataIn2 = 32'd10; 
32'd3306: dataIn2 = 32'd5; 
32'd3307: dataIn2 = 32'd80; 
32'd3308: dataIn2 = 32'd4; 
32'd3309: dataIn2 = 32'd51; 
32'd3310: dataIn2 = 32'd31; 
32'd3311: dataIn2 = 32'd92; 
32'd3312: dataIn2 = 32'd2; 
32'd3313: dataIn2 = 32'd29; 
32'd3314: dataIn2 = 32'd86; 
32'd3315: dataIn2 = 32'd67; 
32'd3316: dataIn2 = 32'd14; 
32'd3317: dataIn2 = 32'd68; 
32'd3318: dataIn2 = 32'd12; 
32'd3319: dataIn2 = 32'd20; 
32'd3320: dataIn2 = 32'd43; 
32'd3321: dataIn2 = 32'd49; 
32'd3322: dataIn2 = 32'd23; 
32'd3323: dataIn2 = 32'd97; 
32'd3324: dataIn2 = 32'd31; 
32'd3325: dataIn2 = 32'd31; 
32'd3326: dataIn2 = 32'd55; 
32'd3327: dataIn2 = 32'd81; 
32'd3328: dataIn2 = 32'd79; 
32'd3329: dataIn2 = 32'd60; 
32'd3330: dataIn2 = 32'd24; 
32'd3331: dataIn2 = 32'd47; 
32'd3332: dataIn2 = 32'd66; 
32'd3333: dataIn2 = 32'd94; 
32'd3334: dataIn2 = 32'd1; 
32'd3335: dataIn2 = 32'd77; 
32'd3336: dataIn2 = 32'd54; 
32'd3337: dataIn2 = 32'd21; 
32'd3338: dataIn2 = 32'd70; 
32'd3339: dataIn2 = 32'd90; 
32'd3340: dataIn2 = 32'd77; 
32'd3341: dataIn2 = 32'd25; 
32'd3342: dataIn2 = 32'd31; 
32'd3343: dataIn2 = 32'd2; 
32'd3344: dataIn2 = 32'd10; 
32'd3345: dataIn2 = 32'd24; 
32'd3346: dataIn2 = 32'd39; 
32'd3347: dataIn2 = 32'd63; 
32'd3348: dataIn2 = 32'd55; 
32'd3349: dataIn2 = 32'd48; 
32'd3350: dataIn2 = 32'd66; 
32'd3351: dataIn2 = 32'd16; 
32'd3352: dataIn2 = 32'd21; 
32'd3353: dataIn2 = 32'd88; 
32'd3354: dataIn2 = 32'd25; 
32'd3355: dataIn2 = 32'd4; 
32'd3356: dataIn2 = 32'd100; 
32'd3357: dataIn2 = 32'd35; 
32'd3358: dataIn2 = 32'd88; 
32'd3359: dataIn2 = 32'd53; 
32'd3360: dataIn2 = 32'd25; 
32'd3361: dataIn2 = 32'd98; 
32'd3362: dataIn2 = 32'd72; 
32'd3363: dataIn2 = 32'd31; 
32'd3364: dataIn2 = 32'd23; 
32'd3365: dataIn2 = 32'd19; 
32'd3366: dataIn2 = 32'd60; 
32'd3367: dataIn2 = 32'd80; 
32'd3368: dataIn2 = 32'd35; 
32'd3369: dataIn2 = 32'd75; 
32'd3370: dataIn2 = 32'd62; 
32'd3371: dataIn2 = 32'd32; 
32'd3372: dataIn2 = 32'd46; 
32'd3373: dataIn2 = 32'd28; 
32'd3374: dataIn2 = 32'd3; 
32'd3375: dataIn2 = 32'd60; 
32'd3376: dataIn2 = 32'd76; 
32'd3377: dataIn2 = 32'd90; 
32'd3378: dataIn2 = 32'd64; 
32'd3379: dataIn2 = 32'd44; 
32'd3380: dataIn2 = 32'd76; 
32'd3381: dataIn2 = 32'd76; 
32'd3382: dataIn2 = 32'd16; 
32'd3383: dataIn2 = 32'd58; 
32'd3384: dataIn2 = 32'd89; 
32'd3385: dataIn2 = 32'd68; 
32'd3386: dataIn2 = 32'd39; 
32'd3387: dataIn2 = 32'd86; 
32'd3388: dataIn2 = 32'd81; 
32'd3389: dataIn2 = 32'd74; 
32'd3390: dataIn2 = 32'd39; 
32'd3391: dataIn2 = 32'd23; 
32'd3392: dataIn2 = 32'd100; 
32'd3393: dataIn2 = 32'd2; 
32'd3394: dataIn2 = 32'd80; 
32'd3395: dataIn2 = 32'd20; 
32'd3396: dataIn2 = 32'd91; 
32'd3397: dataIn2 = 32'd1; 
32'd3398: dataIn2 = 32'd9; 
32'd3399: dataIn2 = 32'd24; 
32'd3400: dataIn2 = 32'd11; 
32'd3401: dataIn2 = 32'd39; 
32'd3402: dataIn2 = 32'd66; 
32'd3403: dataIn2 = 32'd82; 
32'd3404: dataIn2 = 32'd39; 
32'd3405: dataIn2 = 32'd4; 
32'd3406: dataIn2 = 32'd34; 
32'd3407: dataIn2 = 32'd63; 
32'd3408: dataIn2 = 32'd6; 
32'd3409: dataIn2 = 32'd12; 
32'd3410: dataIn2 = 32'd27; 
32'd3411: dataIn2 = 32'd76; 
32'd3412: dataIn2 = 32'd71; 
32'd3413: dataIn2 = 32'd83; 
32'd3414: dataIn2 = 32'd1; 
32'd3415: dataIn2 = 32'd48; 
32'd3416: dataIn2 = 32'd7; 
32'd3417: dataIn2 = 32'd20; 
32'd3418: dataIn2 = 32'd41; 
32'd3419: dataIn2 = 32'd54; 
32'd3420: dataIn2 = 32'd55; 
32'd3421: dataIn2 = 32'd7; 
32'd3422: dataIn2 = 32'd78; 
32'd3423: dataIn2 = 32'd46; 
32'd3424: dataIn2 = 32'd6; 
32'd3425: dataIn2 = 32'd90; 
32'd3426: dataIn2 = 32'd77; 
32'd3427: dataIn2 = 32'd9; 
32'd3428: dataIn2 = 32'd74; 
32'd3429: dataIn2 = 32'd10; 
32'd3430: dataIn2 = 32'd48; 
32'd3431: dataIn2 = 32'd42; 
32'd3432: dataIn2 = 32'd36; 
32'd3433: dataIn2 = 32'd92; 
32'd3434: dataIn2 = 32'd75; 
32'd3435: dataIn2 = 32'd51; 
32'd3436: dataIn2 = 32'd98; 
32'd3437: dataIn2 = 32'd84; 
32'd3438: dataIn2 = 32'd75; 
32'd3439: dataIn2 = 32'd20; 
32'd3440: dataIn2 = 32'd69; 
32'd3441: dataIn2 = 32'd0; 
32'd3442: dataIn2 = 32'd34; 
32'd3443: dataIn2 = 32'd80; 
32'd3444: dataIn2 = 32'd59; 
32'd3445: dataIn2 = 32'd85; 
32'd3446: dataIn2 = 32'd64; 
32'd3447: dataIn2 = 32'd32; 
32'd3448: dataIn2 = 32'd88; 
32'd3449: dataIn2 = 32'd61; 
32'd3450: dataIn2 = 32'd3; 
32'd3451: dataIn2 = 32'd89; 
32'd3452: dataIn2 = 32'd63; 
32'd3453: dataIn2 = 32'd10; 
32'd3454: dataIn2 = 32'd2; 
32'd3455: dataIn2 = 32'd24; 
32'd3456: dataIn2 = 32'd63; 
32'd3457: dataIn2 = 32'd55; 
32'd3458: dataIn2 = 32'd72; 
32'd3459: dataIn2 = 32'd60; 
32'd3460: dataIn2 = 32'd62; 
32'd3461: dataIn2 = 32'd55; 
32'd3462: dataIn2 = 32'd18; 
32'd3463: dataIn2 = 32'd3; 
32'd3464: dataIn2 = 32'd71; 
32'd3465: dataIn2 = 32'd52; 
32'd3466: dataIn2 = 32'd38; 
32'd3467: dataIn2 = 32'd22; 
32'd3468: dataIn2 = 32'd23; 
32'd3469: dataIn2 = 32'd66; 
32'd3470: dataIn2 = 32'd36; 
32'd3471: dataIn2 = 32'd39; 
32'd3472: dataIn2 = 32'd57; 
32'd3473: dataIn2 = 32'd19; 
32'd3474: dataIn2 = 32'd76; 
32'd3475: dataIn2 = 32'd19; 
32'd3476: dataIn2 = 32'd42; 
32'd3477: dataIn2 = 32'd40; 
32'd3478: dataIn2 = 32'd37; 
32'd3479: dataIn2 = 32'd75; 
32'd3480: dataIn2 = 32'd51; 
32'd3481: dataIn2 = 32'd96; 
32'd3482: dataIn2 = 32'd69; 
32'd3483: dataIn2 = 32'd36; 
32'd3484: dataIn2 = 32'd59; 
32'd3485: dataIn2 = 32'd19; 
32'd3486: dataIn2 = 32'd64; 
32'd3487: dataIn2 = 32'd9; 
32'd3488: dataIn2 = 32'd69; 
32'd3489: dataIn2 = 32'd31; 
32'd3490: dataIn2 = 32'd75; 
32'd3491: dataIn2 = 32'd44; 
32'd3492: dataIn2 = 32'd28; 
32'd3493: dataIn2 = 32'd7; 
32'd3494: dataIn2 = 32'd22; 
32'd3495: dataIn2 = 32'd32; 
32'd3496: dataIn2 = 32'd83; 
32'd3497: dataIn2 = 32'd84; 
32'd3498: dataIn2 = 32'd69; 
32'd3499: dataIn2 = 32'd50; 
32'd3500: dataIn2 = 32'd74; 
32'd3501: dataIn2 = 32'd84; 
32'd3502: dataIn2 = 32'd37; 
32'd3503: dataIn2 = 32'd23; 
32'd3504: dataIn2 = 32'd56; 
32'd3505: dataIn2 = 32'd40; 
32'd3506: dataIn2 = 32'd14; 
32'd3507: dataIn2 = 32'd27; 
32'd3508: dataIn2 = 32'd41; 
32'd3509: dataIn2 = 32'd87; 
32'd3510: dataIn2 = 32'd97; 
32'd3511: dataIn2 = 32'd97; 
32'd3512: dataIn2 = 32'd89; 
32'd3513: dataIn2 = 32'd80; 
32'd3514: dataIn2 = 32'd2; 
32'd3515: dataIn2 = 32'd0; 
32'd3516: dataIn2 = 32'd83; 
32'd3517: dataIn2 = 32'd18; 
32'd3518: dataIn2 = 32'd91; 
32'd3519: dataIn2 = 32'd21; 
32'd3520: dataIn2 = 32'd96; 
32'd3521: dataIn2 = 32'd74; 
32'd3522: dataIn2 = 32'd67; 
32'd3523: dataIn2 = 32'd77; 
32'd3524: dataIn2 = 32'd47; 
32'd3525: dataIn2 = 32'd39; 
32'd3526: dataIn2 = 32'd9; 
32'd3527: dataIn2 = 32'd78; 
32'd3528: dataIn2 = 32'd100; 
32'd3529: dataIn2 = 32'd90; 
32'd3530: dataIn2 = 32'd61; 
32'd3531: dataIn2 = 32'd49; 
32'd3532: dataIn2 = 32'd39; 
32'd3533: dataIn2 = 32'd42; 
32'd3534: dataIn2 = 32'd11; 
32'd3535: dataIn2 = 32'd70; 
32'd3536: dataIn2 = 32'd58; 
32'd3537: dataIn2 = 32'd68; 
32'd3538: dataIn2 = 32'd9; 
32'd3539: dataIn2 = 32'd10; 
32'd3540: dataIn2 = 32'd34; 
32'd3541: dataIn2 = 32'd84; 
32'd3542: dataIn2 = 32'd30; 
32'd3543: dataIn2 = 32'd12; 
32'd3544: dataIn2 = 32'd23; 
32'd3545: dataIn2 = 32'd65; 
32'd3546: dataIn2 = 32'd33; 
32'd3547: dataIn2 = 32'd14; 
32'd3548: dataIn2 = 32'd1; 
32'd3549: dataIn2 = 32'd9; 
32'd3550: dataIn2 = 32'd57; 
32'd3551: dataIn2 = 32'd76; 
32'd3552: dataIn2 = 32'd44; 
32'd3553: dataIn2 = 32'd98; 
32'd3554: dataIn2 = 32'd22; 
32'd3555: dataIn2 = 32'd51; 
32'd3556: dataIn2 = 32'd48; 
32'd3557: dataIn2 = 32'd74; 
32'd3558: dataIn2 = 32'd39; 
32'd3559: dataIn2 = 32'd63; 
32'd3560: dataIn2 = 32'd28; 
32'd3561: dataIn2 = 32'd49; 
32'd3562: dataIn2 = 32'd44; 
32'd3563: dataIn2 = 32'd98; 
32'd3564: dataIn2 = 32'd71; 
32'd3565: dataIn2 = 32'd10; 
32'd3566: dataIn2 = 32'd2; 
32'd3567: dataIn2 = 32'd66; 
32'd3568: dataIn2 = 32'd50; 
32'd3569: dataIn2 = 32'd100; 
32'd3570: dataIn2 = 32'd10; 
32'd3571: dataIn2 = 32'd89; 
32'd3572: dataIn2 = 32'd66; 
32'd3573: dataIn2 = 32'd31; 
32'd3574: dataIn2 = 32'd51; 
32'd3575: dataIn2 = 32'd50; 
32'd3576: dataIn2 = 32'd89; 
32'd3577: dataIn2 = 32'd68; 
32'd3578: dataIn2 = 32'd41; 
32'd3579: dataIn2 = 32'd5; 
32'd3580: dataIn2 = 32'd63; 
32'd3581: dataIn2 = 32'd78; 
32'd3582: dataIn2 = 32'd16; 
32'd3583: dataIn2 = 32'd8; 
32'd3584: dataIn2 = 32'd77; 
32'd3585: dataIn2 = 32'd93; 
32'd3586: dataIn2 = 32'd98; 
32'd3587: dataIn2 = 32'd25; 
32'd3588: dataIn2 = 32'd2; 
32'd3589: dataIn2 = 32'd18; 
32'd3590: dataIn2 = 32'd33; 
32'd3591: dataIn2 = 32'd75; 
32'd3592: dataIn2 = 32'd93; 
32'd3593: dataIn2 = 32'd79; 
32'd3594: dataIn2 = 32'd84; 
32'd3595: dataIn2 = 32'd54; 
32'd3596: dataIn2 = 32'd92; 
32'd3597: dataIn2 = 32'd6; 
32'd3598: dataIn2 = 32'd97; 
32'd3599: dataIn2 = 32'd55; 
32'd3600: dataIn2 = 32'd98; 
32'd3601: dataIn2 = 32'd55; 
32'd3602: dataIn2 = 32'd16; 
32'd3603: dataIn2 = 32'd35; 
32'd3604: dataIn2 = 32'd74; 
32'd3605: dataIn2 = 32'd29; 
32'd3606: dataIn2 = 32'd30; 
32'd3607: dataIn2 = 32'd55; 
32'd3608: dataIn2 = 32'd49; 
32'd3609: dataIn2 = 32'd86; 
32'd3610: dataIn2 = 32'd73; 
32'd3611: dataIn2 = 32'd21; 
32'd3612: dataIn2 = 32'd98; 
32'd3613: dataIn2 = 32'd6; 
32'd3614: dataIn2 = 32'd63; 
32'd3615: dataIn2 = 32'd27; 
32'd3616: dataIn2 = 32'd6; 
32'd3617: dataIn2 = 32'd45; 
32'd3618: dataIn2 = 32'd75; 
32'd3619: dataIn2 = 32'd50; 
32'd3620: dataIn2 = 32'd32; 
32'd3621: dataIn2 = 32'd20; 
32'd3622: dataIn2 = 32'd60; 
32'd3623: dataIn2 = 32'd38; 
32'd3624: dataIn2 = 32'd60; 
32'd3625: dataIn2 = 32'd57; 
32'd3626: dataIn2 = 32'd38; 
32'd3627: dataIn2 = 32'd92; 
32'd3628: dataIn2 = 32'd34; 
32'd3629: dataIn2 = 32'd83; 
32'd3630: dataIn2 = 32'd10; 
32'd3631: dataIn2 = 32'd10; 
32'd3632: dataIn2 = 32'd2; 
32'd3633: dataIn2 = 32'd60; 
32'd3634: dataIn2 = 32'd17; 
32'd3635: dataIn2 = 32'd65; 
32'd3636: dataIn2 = 32'd16; 
32'd3637: dataIn2 = 32'd51; 
32'd3638: dataIn2 = 32'd79; 
32'd3639: dataIn2 = 32'd7; 
32'd3640: dataIn2 = 32'd98; 
32'd3641: dataIn2 = 32'd58; 
32'd3642: dataIn2 = 32'd76; 
32'd3643: dataIn2 = 32'd81; 
32'd3644: dataIn2 = 32'd84; 
32'd3645: dataIn2 = 32'd46; 
32'd3646: dataIn2 = 32'd20; 
32'd3647: dataIn2 = 32'd92; 
32'd3648: dataIn2 = 32'd15; 
32'd3649: dataIn2 = 32'd23; 
32'd3650: dataIn2 = 32'd37; 
32'd3651: dataIn2 = 32'd78; 
32'd3652: dataIn2 = 32'd31; 
32'd3653: dataIn2 = 32'd72; 
32'd3654: dataIn2 = 32'd72; 
32'd3655: dataIn2 = 32'd58; 
32'd3656: dataIn2 = 32'd52; 
32'd3657: dataIn2 = 32'd72; 
32'd3658: dataIn2 = 32'd90; 
32'd3659: dataIn2 = 32'd90; 
32'd3660: dataIn2 = 32'd12; 
32'd3661: dataIn2 = 32'd35; 
32'd3662: dataIn2 = 32'd59; 
32'd3663: dataIn2 = 32'd72; 
32'd3664: dataIn2 = 32'd71; 
32'd3665: dataIn2 = 32'd84; 
32'd3666: dataIn2 = 32'd79; 
32'd3667: dataIn2 = 32'd10; 
32'd3668: dataIn2 = 32'd100; 
32'd3669: dataIn2 = 32'd47; 
32'd3670: dataIn2 = 32'd17; 
32'd3671: dataIn2 = 32'd26; 
32'd3672: dataIn2 = 32'd72; 
32'd3673: dataIn2 = 32'd96; 
32'd3674: dataIn2 = 32'd63; 
32'd3675: dataIn2 = 32'd12; 
32'd3676: dataIn2 = 32'd97; 
32'd3677: dataIn2 = 32'd22; 
32'd3678: dataIn2 = 32'd30; 
32'd3679: dataIn2 = 32'd15; 
32'd3680: dataIn2 = 32'd96; 
32'd3681: dataIn2 = 32'd15; 
32'd3682: dataIn2 = 32'd0; 
32'd3683: dataIn2 = 32'd27; 
32'd3684: dataIn2 = 32'd70; 
32'd3685: dataIn2 = 32'd79; 
32'd3686: dataIn2 = 32'd67; 
32'd3687: dataIn2 = 32'd22; 
32'd3688: dataIn2 = 32'd18; 
32'd3689: dataIn2 = 32'd30; 
32'd3690: dataIn2 = 32'd70; 
32'd3691: dataIn2 = 32'd97; 
32'd3692: dataIn2 = 32'd99; 
32'd3693: dataIn2 = 32'd97; 
32'd3694: dataIn2 = 32'd50; 
32'd3695: dataIn2 = 32'd43; 
32'd3696: dataIn2 = 32'd39; 
32'd3697: dataIn2 = 32'd70; 
32'd3698: dataIn2 = 32'd15; 
32'd3699: dataIn2 = 32'd88; 
32'd3700: dataIn2 = 32'd55; 
32'd3701: dataIn2 = 32'd24; 
32'd3702: dataIn2 = 32'd86; 
32'd3703: dataIn2 = 32'd32; 
32'd3704: dataIn2 = 32'd38; 
32'd3705: dataIn2 = 32'd21; 
32'd3706: dataIn2 = 32'd92; 
32'd3707: dataIn2 = 32'd24; 
32'd3708: dataIn2 = 32'd34; 
32'd3709: dataIn2 = 32'd64; 
32'd3710: dataIn2 = 32'd48; 
32'd3711: dataIn2 = 32'd8; 
32'd3712: dataIn2 = 32'd69; 
32'd3713: dataIn2 = 32'd98; 
32'd3714: dataIn2 = 32'd31; 
32'd3715: dataIn2 = 32'd73; 
32'd3716: dataIn2 = 32'd45; 
32'd3717: dataIn2 = 32'd34; 
32'd3718: dataIn2 = 32'd73; 
32'd3719: dataIn2 = 32'd85; 
32'd3720: dataIn2 = 32'd29; 
32'd3721: dataIn2 = 32'd14; 
32'd3722: dataIn2 = 32'd7; 
32'd3723: dataIn2 = 32'd36; 
32'd3724: dataIn2 = 32'd76; 
32'd3725: dataIn2 = 32'd59; 
32'd3726: dataIn2 = 32'd30; 
32'd3727: dataIn2 = 32'd42; 
32'd3728: dataIn2 = 32'd19; 
32'd3729: dataIn2 = 32'd39; 
32'd3730: dataIn2 = 32'd49; 
32'd3731: dataIn2 = 32'd44; 
32'd3732: dataIn2 = 32'd37; 
32'd3733: dataIn2 = 32'd60; 
32'd3734: dataIn2 = 32'd67; 
32'd3735: dataIn2 = 32'd91; 
32'd3736: dataIn2 = 32'd78; 
32'd3737: dataIn2 = 32'd61; 
32'd3738: dataIn2 = 32'd43; 
32'd3739: dataIn2 = 32'd73; 
32'd3740: dataIn2 = 32'd86; 
32'd3741: dataIn2 = 32'd81; 
32'd3742: dataIn2 = 32'd57; 
32'd3743: dataIn2 = 32'd84; 
32'd3744: dataIn2 = 32'd83; 
32'd3745: dataIn2 = 32'd46; 
32'd3746: dataIn2 = 32'd65; 
32'd3747: dataIn2 = 32'd73; 
32'd3748: dataIn2 = 32'd18; 
32'd3749: dataIn2 = 32'd74; 
32'd3750: dataIn2 = 32'd31; 
32'd3751: dataIn2 = 32'd45; 
32'd3752: dataIn2 = 32'd41; 
32'd3753: dataIn2 = 32'd88; 
32'd3754: dataIn2 = 32'd35; 
32'd3755: dataIn2 = 32'd49; 
32'd3756: dataIn2 = 32'd90; 
32'd3757: dataIn2 = 32'd40; 
32'd3758: dataIn2 = 32'd0; 
32'd3759: dataIn2 = 32'd7; 
32'd3760: dataIn2 = 32'd97; 
32'd3761: dataIn2 = 32'd85; 
32'd3762: dataIn2 = 32'd49; 
32'd3763: dataIn2 = 32'd20; 
32'd3764: dataIn2 = 32'd46; 
32'd3765: dataIn2 = 32'd13; 
32'd3766: dataIn2 = 32'd20; 
32'd3767: dataIn2 = 32'd20; 
32'd3768: dataIn2 = 32'd80; 
32'd3769: dataIn2 = 32'd40; 
32'd3770: dataIn2 = 32'd89; 
32'd3771: dataIn2 = 32'd9; 
32'd3772: dataIn2 = 32'd51; 
32'd3773: dataIn2 = 32'd63; 
32'd3774: dataIn2 = 32'd49; 
32'd3775: dataIn2 = 32'd17; 
32'd3776: dataIn2 = 32'd54; 
32'd3777: dataIn2 = 32'd30; 
32'd3778: dataIn2 = 32'd22; 
32'd3779: dataIn2 = 32'd0; 
32'd3780: dataIn2 = 32'd7; 
32'd3781: dataIn2 = 32'd20; 
32'd3782: dataIn2 = 32'd24; 
32'd3783: dataIn2 = 32'd72; 
32'd3784: dataIn2 = 32'd19; 
32'd3785: dataIn2 = 32'd16; 
32'd3786: dataIn2 = 32'd78; 
32'd3787: dataIn2 = 32'd80; 
32'd3788: dataIn2 = 32'd28; 
32'd3789: dataIn2 = 32'd60; 
32'd3790: dataIn2 = 32'd6; 
32'd3791: dataIn2 = 32'd20; 
32'd3792: dataIn2 = 32'd74; 
32'd3793: dataIn2 = 32'd61; 
32'd3794: dataIn2 = 32'd10; 
32'd3795: dataIn2 = 32'd74; 
32'd3796: dataIn2 = 32'd66; 
32'd3797: dataIn2 = 32'd22; 
32'd3798: dataIn2 = 32'd83; 
32'd3799: dataIn2 = 32'd66; 
32'd3800: dataIn2 = 32'd84; 
32'd3801: dataIn2 = 32'd18; 
32'd3802: dataIn2 = 32'd79; 
32'd3803: dataIn2 = 32'd67; 
32'd3804: dataIn2 = 32'd31; 
32'd3805: dataIn2 = 32'd18; 
32'd3806: dataIn2 = 32'd28; 
32'd3807: dataIn2 = 32'd76; 
32'd3808: dataIn2 = 32'd79; 
32'd3809: dataIn2 = 32'd74; 
32'd3810: dataIn2 = 32'd17; 
32'd3811: dataIn2 = 32'd29; 
32'd3812: dataIn2 = 32'd57; 
32'd3813: dataIn2 = 32'd4; 
32'd3814: dataIn2 = 32'd21; 
32'd3815: dataIn2 = 32'd71; 
32'd3816: dataIn2 = 32'd79; 
32'd3817: dataIn2 = 32'd55; 
32'd3818: dataIn2 = 32'd65; 
32'd3819: dataIn2 = 32'd7; 
32'd3820: dataIn2 = 32'd40; 
32'd3821: dataIn2 = 32'd13; 
32'd3822: dataIn2 = 32'd27; 
32'd3823: dataIn2 = 32'd60; 
32'd3824: dataIn2 = 32'd95; 
32'd3825: dataIn2 = 32'd70; 
32'd3826: dataIn2 = 32'd77; 
32'd3827: dataIn2 = 32'd75; 
32'd3828: dataIn2 = 32'd17; 
32'd3829: dataIn2 = 32'd62; 
32'd3830: dataIn2 = 32'd44; 
32'd3831: dataIn2 = 32'd61; 
32'd3832: dataIn2 = 32'd21; 
32'd3833: dataIn2 = 32'd66; 
32'd3834: dataIn2 = 32'd25; 
32'd3835: dataIn2 = 32'd31; 
32'd3836: dataIn2 = 32'd76; 
32'd3837: dataIn2 = 32'd99; 
32'd3838: dataIn2 = 32'd13; 
32'd3839: dataIn2 = 32'd29; 
32'd3840: dataIn2 = 32'd53; 
32'd3841: dataIn2 = 32'd48; 
32'd3842: dataIn2 = 32'd53; 
32'd3843: dataIn2 = 32'd9; 
32'd3844: dataIn2 = 32'd52; 
32'd3845: dataIn2 = 32'd83; 
32'd3846: dataIn2 = 32'd55; 
32'd3847: dataIn2 = 32'd14; 
32'd3848: dataIn2 = 32'd23; 
32'd3849: dataIn2 = 32'd97; 
32'd3850: dataIn2 = 32'd1; 
32'd3851: dataIn2 = 32'd54; 
32'd3852: dataIn2 = 32'd5; 
32'd3853: dataIn2 = 32'd7; 
32'd3854: dataIn2 = 32'd86; 
32'd3855: dataIn2 = 32'd91; 
32'd3856: dataIn2 = 32'd66; 
32'd3857: dataIn2 = 32'd64; 
32'd3858: dataIn2 = 32'd68; 
32'd3859: dataIn2 = 32'd23; 
32'd3860: dataIn2 = 32'd14; 
32'd3861: dataIn2 = 32'd68; 
32'd3862: dataIn2 = 32'd50; 
32'd3863: dataIn2 = 32'd19; 
32'd3864: dataIn2 = 32'd75; 
32'd3865: dataIn2 = 32'd89; 
32'd3866: dataIn2 = 32'd52; 
32'd3867: dataIn2 = 32'd64; 
32'd3868: dataIn2 = 32'd35; 
32'd3869: dataIn2 = 32'd62; 
32'd3870: dataIn2 = 32'd0; 
32'd3871: dataIn2 = 32'd33; 
32'd3872: dataIn2 = 32'd81; 
32'd3873: dataIn2 = 32'd41; 
32'd3874: dataIn2 = 32'd86; 
32'd3875: dataIn2 = 32'd19; 
32'd3876: dataIn2 = 32'd98; 
32'd3877: dataIn2 = 32'd29; 
32'd3878: dataIn2 = 32'd17; 
32'd3879: dataIn2 = 32'd88; 
32'd3880: dataIn2 = 32'd88; 
32'd3881: dataIn2 = 32'd79; 
32'd3882: dataIn2 = 32'd52; 
32'd3883: dataIn2 = 32'd51; 
32'd3884: dataIn2 = 32'd46; 
32'd3885: dataIn2 = 32'd60; 
32'd3886: dataIn2 = 32'd45; 
32'd3887: dataIn2 = 32'd12; 
32'd3888: dataIn2 = 32'd59; 
32'd3889: dataIn2 = 32'd94; 
32'd3890: dataIn2 = 32'd34; 
32'd3891: dataIn2 = 32'd16; 
32'd3892: dataIn2 = 32'd20; 
32'd3893: dataIn2 = 32'd12; 
32'd3894: dataIn2 = 32'd45; 
32'd3895: dataIn2 = 32'd75; 
32'd3896: dataIn2 = 32'd0; 
32'd3897: dataIn2 = 32'd55; 
32'd3898: dataIn2 = 32'd81; 
32'd3899: dataIn2 = 32'd10; 
32'd3900: dataIn2 = 32'd65; 
32'd3901: dataIn2 = 32'd71; 
32'd3902: dataIn2 = 32'd12; 
32'd3903: dataIn2 = 32'd10; 
32'd3904: dataIn2 = 32'd83; 
32'd3905: dataIn2 = 32'd55; 
32'd3906: dataIn2 = 32'd67; 
32'd3907: dataIn2 = 32'd45; 
32'd3908: dataIn2 = 32'd31; 
32'd3909: dataIn2 = 32'd58; 
32'd3910: dataIn2 = 32'd25; 
32'd3911: dataIn2 = 32'd28; 
32'd3912: dataIn2 = 32'd65; 
32'd3913: dataIn2 = 32'd11; 
32'd3914: dataIn2 = 32'd84; 
32'd3915: dataIn2 = 32'd65; 
32'd3916: dataIn2 = 32'd48; 
32'd3917: dataIn2 = 32'd51; 
32'd3918: dataIn2 = 32'd81; 
32'd3919: dataIn2 = 32'd91; 
32'd3920: dataIn2 = 32'd58; 
32'd3921: dataIn2 = 32'd58; 
32'd3922: dataIn2 = 32'd81; 
32'd3923: dataIn2 = 32'd50; 
32'd3924: dataIn2 = 32'd97; 
32'd3925: dataIn2 = 32'd69; 
32'd3926: dataIn2 = 32'd28; 
32'd3927: dataIn2 = 32'd38; 
32'd3928: dataIn2 = 32'd34; 
32'd3929: dataIn2 = 32'd97; 
32'd3930: dataIn2 = 32'd62; 
32'd3931: dataIn2 = 32'd13; 
32'd3932: dataIn2 = 32'd27; 
32'd3933: dataIn2 = 32'd1; 
32'd3934: dataIn2 = 32'd33; 
32'd3935: dataIn2 = 32'd13; 
32'd3936: dataIn2 = 32'd43; 
32'd3937: dataIn2 = 32'd83; 
32'd3938: dataIn2 = 32'd44; 
32'd3939: dataIn2 = 32'd95; 
32'd3940: dataIn2 = 32'd59; 
32'd3941: dataIn2 = 32'd78; 
32'd3942: dataIn2 = 32'd24; 
32'd3943: dataIn2 = 32'd9; 
32'd3944: dataIn2 = 32'd55; 
32'd3945: dataIn2 = 32'd69; 
32'd3946: dataIn2 = 32'd73; 
32'd3947: dataIn2 = 32'd19; 
32'd3948: dataIn2 = 32'd11; 
32'd3949: dataIn2 = 32'd99; 
32'd3950: dataIn2 = 32'd27; 
32'd3951: dataIn2 = 32'd21; 
32'd3952: dataIn2 = 32'd39; 
32'd3953: dataIn2 = 32'd34; 
32'd3954: dataIn2 = 32'd14; 
32'd3955: dataIn2 = 32'd54; 
32'd3956: dataIn2 = 32'd63; 
32'd3957: dataIn2 = 32'd10; 
32'd3958: dataIn2 = 32'd55; 
32'd3959: dataIn2 = 32'd14; 
32'd3960: dataIn2 = 32'd0; 
32'd3961: dataIn2 = 32'd81; 
32'd3962: dataIn2 = 32'd60; 
32'd3963: dataIn2 = 32'd32; 
32'd3964: dataIn2 = 32'd76; 
32'd3965: dataIn2 = 32'd75; 
32'd3966: dataIn2 = 32'd19; 
32'd3967: dataIn2 = 32'd70; 
32'd3968: dataIn2 = 32'd23; 
32'd3969: dataIn2 = 32'd5; 
32'd3970: dataIn2 = 32'd52; 
32'd3971: dataIn2 = 32'd93; 
32'd3972: dataIn2 = 32'd39; 
32'd3973: dataIn2 = 32'd78; 
32'd3974: dataIn2 = 32'd67; 
32'd3975: dataIn2 = 32'd47; 
32'd3976: dataIn2 = 32'd66; 
32'd3977: dataIn2 = 32'd42; 
32'd3978: dataIn2 = 32'd18; 
32'd3979: dataIn2 = 32'd49; 
32'd3980: dataIn2 = 32'd12; 
32'd3981: dataIn2 = 32'd39; 
32'd3982: dataIn2 = 32'd13; 
32'd3983: dataIn2 = 32'd59; 
32'd3984: dataIn2 = 32'd7; 
32'd3985: dataIn2 = 32'd74; 
32'd3986: dataIn2 = 32'd68; 
32'd3987: dataIn2 = 32'd24; 
32'd3988: dataIn2 = 32'd24; 
32'd3989: dataIn2 = 32'd0; 
32'd3990: dataIn2 = 32'd85; 
32'd3991: dataIn2 = 32'd21; 
32'd3992: dataIn2 = 32'd3; 
32'd3993: dataIn2 = 32'd8; 
32'd3994: dataIn2 = 32'd64; 
32'd3995: dataIn2 = 32'd59; 
32'd3996: dataIn2 = 32'd60; 
32'd3997: dataIn2 = 32'd33; 
32'd3998: dataIn2 = 32'd53; 
32'd3999: dataIn2 = 32'd98; 
32'd4000: dataIn2 = 32'd72; 
32'd4001: dataIn2 = 32'd9; 
32'd4002: dataIn2 = 32'd5; 
32'd4003: dataIn2 = 32'd4; 
32'd4004: dataIn2 = 32'd36; 
32'd4005: dataIn2 = 32'd6; 
32'd4006: dataIn2 = 32'd21; 
32'd4007: dataIn2 = 32'd80; 
32'd4008: dataIn2 = 32'd8; 
32'd4009: dataIn2 = 32'd95; 
32'd4010: dataIn2 = 32'd91; 
32'd4011: dataIn2 = 32'd80; 
32'd4012: dataIn2 = 32'd53; 
32'd4013: dataIn2 = 32'd64; 
32'd4014: dataIn2 = 32'd67; 
32'd4015: dataIn2 = 32'd24; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_64_10.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
