//64x64 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 819 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd330 ; 
  wdata_col_base = 32'd11490 ; 
  row_base = 32'd123090 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #96800; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd123090: dataIn1 = 32'd0
; 
32'd123091: dataIn1 = 32'd14
; 
32'd123092: dataIn1 = 32'd27
; 
32'd123093: dataIn1 = 32'd43
; 
32'd123094: dataIn1 = 32'd51
; 
32'd123095: dataIn1 = 32'd64
; 
32'd123096: dataIn1 = 32'd74
; 
32'd123097: dataIn1 = 32'd83
; 
32'd123098: dataIn1 = 32'd97
; 
32'd123099: dataIn1 = 32'd108
; 
32'd123100: dataIn1 = 32'd124
; 
32'd123101: dataIn1 = 32'd134
; 
32'd123102: dataIn1 = 32'd142
; 
32'd123103: dataIn1 = 32'd155
; 
32'd123104: dataIn1 = 32'd169
; 
32'd123105: dataIn1 = 32'd178
; 
32'd123106: dataIn1 = 32'd194
; 
32'd123107: dataIn1 = 32'd212
; 
32'd123108: dataIn1 = 32'd221
; 
32'd123109: dataIn1 = 32'd236
; 
32'd123110: dataIn1 = 32'd246
; 
32'd123111: dataIn1 = 32'd257
; 
32'd123112: dataIn1 = 32'd271
; 
32'd123113: dataIn1 = 32'd287
; 
32'd123114: dataIn1 = 32'd302
; 
32'd123115: dataIn1 = 32'd317
; 
32'd123116: dataIn1 = 32'd333
; 
32'd123117: dataIn1 = 32'd351
; 
32'd123118: dataIn1 = 32'd361
; 
32'd123119: dataIn1 = 32'd370
; 
32'd123120: dataIn1 = 32'd380
; 
32'd123121: dataIn1 = 32'd391
; 
32'd123122: dataIn1 = 32'd400
; 
32'd123123: dataIn1 = 32'd413
; 
32'd123124: dataIn1 = 32'd432
; 
32'd123125: dataIn1 = 32'd445
; 
32'd123126: dataIn1 = 32'd458
; 
32'd123127: dataIn1 = 32'd472
; 
32'd123128: dataIn1 = 32'd483
; 
32'd123129: dataIn1 = 32'd495
; 
32'd123130: dataIn1 = 32'd504
; 
32'd123131: dataIn1 = 32'd521
; 
32'd123132: dataIn1 = 32'd533
; 
32'd123133: dataIn1 = 32'd544
; 
32'd123134: dataIn1 = 32'd553
; 
32'd123135: dataIn1 = 32'd566
; 
32'd123136: dataIn1 = 32'd580
; 
32'd123137: dataIn1 = 32'd593
; 
32'd123138: dataIn1 = 32'd607
; 
32'd123139: dataIn1 = 32'd616
; 
32'd123140: dataIn1 = 32'd626
; 
32'd123141: dataIn1 = 32'd639
; 
32'd123142: dataIn1 = 32'd652
; 
32'd123143: dataIn1 = 32'd671
; 
32'd123144: dataIn1 = 32'd687
; 
32'd123145: dataIn1 = 32'd699
; 
32'd123146: dataIn1 = 32'd710
; 
32'd123147: dataIn1 = 32'd721
; 
32'd123148: dataIn1 = 32'd734
; 
32'd123149: dataIn1 = 32'd747
; 
32'd123150: dataIn1 = 32'd757
; 
32'd123151: dataIn1 = 32'd767
; 
32'd123152: dataIn1 = 32'd785
; 
32'd123153: dataIn1 = 32'd797
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd11490: dataIn1 = 32'd0
; 
32'd11491: dataIn1 = 32'd14
; 
32'd11492: dataIn1 = 32'd27
; 
32'd11493: dataIn1 = 32'd43
; 
32'd11494: dataIn1 = 32'd51
; 
32'd11495: dataIn1 = 32'd64
; 
32'd11496: dataIn1 = 32'd74
; 
32'd11497: dataIn1 = 32'd83
; 
32'd11498: dataIn1 = 32'd97
; 
32'd11499: dataIn1 = 32'd108
; 
32'd11500: dataIn1 = 32'd124
; 
32'd11501: dataIn1 = 32'd134
; 
32'd11502: dataIn1 = 32'd142
; 
32'd11503: dataIn1 = 32'd155
; 
32'd11504: dataIn1 = 32'd169
; 
32'd11505: dataIn1 = 32'd178
; 
32'd11506: dataIn1 = 32'd194
; 
32'd11507: dataIn1 = 32'd212
; 
32'd11508: dataIn1 = 32'd221
; 
32'd11509: dataIn1 = 32'd236
; 
32'd11510: dataIn1 = 32'd246
; 
32'd11511: dataIn1 = 32'd257
; 
32'd11512: dataIn1 = 32'd271
; 
32'd11513: dataIn1 = 32'd287
; 
32'd11514: dataIn1 = 32'd302
; 
32'd11515: dataIn1 = 32'd317
; 
32'd11516: dataIn1 = 32'd333
; 
32'd11517: dataIn1 = 32'd351
; 
32'd11518: dataIn1 = 32'd361
; 
32'd11519: dataIn1 = 32'd370
; 
32'd11520: dataIn1 = 32'd380
; 
32'd11521: dataIn1 = 32'd391
; 
32'd11522: dataIn1 = 32'd400
; 
32'd11523: dataIn1 = 32'd413
; 
32'd11524: dataIn1 = 32'd432
; 
32'd11525: dataIn1 = 32'd445
; 
32'd11526: dataIn1 = 32'd458
; 
32'd11527: dataIn1 = 32'd472
; 
32'd11528: dataIn1 = 32'd483
; 
32'd11529: dataIn1 = 32'd495
; 
32'd11530: dataIn1 = 32'd504
; 
32'd11531: dataIn1 = 32'd521
; 
32'd11532: dataIn1 = 32'd533
; 
32'd11533: dataIn1 = 32'd544
; 
32'd11534: dataIn1 = 32'd553
; 
32'd11535: dataIn1 = 32'd566
; 
32'd11536: dataIn1 = 32'd580
; 
32'd11537: dataIn1 = 32'd593
; 
32'd11538: dataIn1 = 32'd607
; 
32'd11539: dataIn1 = 32'd616
; 
32'd11540: dataIn1 = 32'd626
; 
32'd11541: dataIn1 = 32'd639
; 
32'd11542: dataIn1 = 32'd652
; 
32'd11543: dataIn1 = 32'd671
; 
32'd11544: dataIn1 = 32'd687
; 
32'd11545: dataIn1 = 32'd699
; 
32'd11546: dataIn1 = 32'd710
; 
32'd11547: dataIn1 = 32'd721
; 
32'd11548: dataIn1 = 32'd734
; 
32'd11549: dataIn1 = 32'd747
; 
32'd11550: dataIn1 = 32'd757
; 
32'd11551: dataIn1 = 32'd767
; 
32'd11552: dataIn1 = 32'd785
; 
32'd11553: dataIn1 = 32'd797
; 
32'd11554: dataIn1 = 32'd812
; 
32'd11555: dataIn1 = 32'd4
; 
32'd11556: dataIn1 = 32'd7
; 
32'd11557: dataIn1 = 32'd8
; 
32'd11558: dataIn1 = 32'd27
; 
32'd11559: dataIn1 = 32'd33
; 
32'd11560: dataIn1 = 32'd44
; 
32'd11561: dataIn1 = 32'd45
; 
32'd11562: dataIn1 = 32'd49
; 
32'd11563: dataIn1 = 32'd51
; 
32'd11564: dataIn1 = 32'd52
; 
32'd11565: dataIn1 = 32'd54
; 
32'd11566: dataIn1 = 32'd55
; 
32'd11567: dataIn1 = 32'd62
; 
32'd11568: dataIn1 = 32'd63
; 
32'd11569: dataIn1 = 32'd0
; 
32'd11570: dataIn1 = 32'd11
; 
32'd11571: dataIn1 = 32'd12
; 
32'd11572: dataIn1 = 32'd21
; 
32'd11573: dataIn1 = 32'd29
; 
32'd11574: dataIn1 = 32'd31
; 
32'd11575: dataIn1 = 32'd40
; 
32'd11576: dataIn1 = 32'd43
; 
32'd11577: dataIn1 = 32'd45
; 
32'd11578: dataIn1 = 32'd56
; 
32'd11579: dataIn1 = 32'd57
; 
32'd11580: dataIn1 = 32'd58
; 
32'd11581: dataIn1 = 32'd60
; 
32'd11582: dataIn1 = 32'd1
; 
32'd11583: dataIn1 = 32'd4
; 
32'd11584: dataIn1 = 32'd7
; 
32'd11585: dataIn1 = 32'd11
; 
32'd11586: dataIn1 = 32'd12
; 
32'd11587: dataIn1 = 32'd14
; 
32'd11588: dataIn1 = 32'd19
; 
32'd11589: dataIn1 = 32'd21
; 
32'd11590: dataIn1 = 32'd24
; 
32'd11591: dataIn1 = 32'd29
; 
32'd11592: dataIn1 = 32'd32
; 
32'd11593: dataIn1 = 32'd34
; 
32'd11594: dataIn1 = 32'd54
; 
32'd11595: dataIn1 = 32'd59
; 
32'd11596: dataIn1 = 32'd61
; 
32'd11597: dataIn1 = 32'd62
; 
32'd11598: dataIn1 = 32'd3
; 
32'd11599: dataIn1 = 32'd9
; 
32'd11600: dataIn1 = 32'd10
; 
32'd11601: dataIn1 = 32'd17
; 
32'd11602: dataIn1 = 32'd29
; 
32'd11603: dataIn1 = 32'd31
; 
32'd11604: dataIn1 = 32'd52
; 
32'd11605: dataIn1 = 32'd55
; 
32'd11606: dataIn1 = 32'd1
; 
32'd11607: dataIn1 = 32'd7
; 
32'd11608: dataIn1 = 32'd10
; 
32'd11609: dataIn1 = 32'd16
; 
32'd11610: dataIn1 = 32'd17
; 
32'd11611: dataIn1 = 32'd18
; 
32'd11612: dataIn1 = 32'd21
; 
32'd11613: dataIn1 = 32'd40
; 
32'd11614: dataIn1 = 32'd42
; 
32'd11615: dataIn1 = 32'd44
; 
32'd11616: dataIn1 = 32'd50
; 
32'd11617: dataIn1 = 32'd54
; 
32'd11618: dataIn1 = 32'd58
; 
32'd11619: dataIn1 = 32'd4
; 
32'd11620: dataIn1 = 32'd11
; 
32'd11621: dataIn1 = 32'd12
; 
32'd11622: dataIn1 = 32'd13
; 
32'd11623: dataIn1 = 32'd42
; 
32'd11624: dataIn1 = 32'd56
; 
32'd11625: dataIn1 = 32'd57
; 
32'd11626: dataIn1 = 32'd60
; 
32'd11627: dataIn1 = 32'd61
; 
32'd11628: dataIn1 = 32'd62
; 
32'd11629: dataIn1 = 32'd2
; 
32'd11630: dataIn1 = 32'd6
; 
32'd11631: dataIn1 = 32'd11
; 
32'd11632: dataIn1 = 32'd12
; 
32'd11633: dataIn1 = 32'd14
; 
32'd11634: dataIn1 = 32'd16
; 
32'd11635: dataIn1 = 32'd27
; 
32'd11636: dataIn1 = 32'd37
; 
32'd11637: dataIn1 = 32'd46
; 
32'd11638: dataIn1 = 32'd4
; 
32'd11639: dataIn1 = 32'd10
; 
32'd11640: dataIn1 = 32'd14
; 
32'd11641: dataIn1 = 32'd16
; 
32'd11642: dataIn1 = 32'd17
; 
32'd11643: dataIn1 = 32'd19
; 
32'd11644: dataIn1 = 32'd37
; 
32'd11645: dataIn1 = 32'd44
; 
32'd11646: dataIn1 = 32'd47
; 
32'd11647: dataIn1 = 32'd48
; 
32'd11648: dataIn1 = 32'd49
; 
32'd11649: dataIn1 = 32'd50
; 
32'd11650: dataIn1 = 32'd53
; 
32'd11651: dataIn1 = 32'd54
; 
32'd11652: dataIn1 = 32'd6
; 
32'd11653: dataIn1 = 32'd14
; 
32'd11654: dataIn1 = 32'd23
; 
32'd11655: dataIn1 = 32'd27
; 
32'd11656: dataIn1 = 32'd29
; 
32'd11657: dataIn1 = 32'd33
; 
32'd11658: dataIn1 = 32'd43
; 
32'd11659: dataIn1 = 32'd44
; 
32'd11660: dataIn1 = 32'd45
; 
32'd11661: dataIn1 = 32'd56
; 
32'd11662: dataIn1 = 32'd63
; 
32'd11663: dataIn1 = 32'd2
; 
32'd11664: dataIn1 = 32'd5
; 
32'd11665: dataIn1 = 32'd9
; 
32'd11666: dataIn1 = 32'd12
; 
32'd11667: dataIn1 = 32'd14
; 
32'd11668: dataIn1 = 32'd20
; 
32'd11669: dataIn1 = 32'd21
; 
32'd11670: dataIn1 = 32'd24
; 
32'd11671: dataIn1 = 32'd29
; 
32'd11672: dataIn1 = 32'd31
; 
32'd11673: dataIn1 = 32'd35
; 
32'd11674: dataIn1 = 32'd44
; 
32'd11675: dataIn1 = 32'd52
; 
32'd11676: dataIn1 = 32'd54
; 
32'd11677: dataIn1 = 32'd58
; 
32'd11678: dataIn1 = 32'd59
; 
32'd11679: dataIn1 = 32'd2
; 
32'd11680: dataIn1 = 32'd3
; 
32'd11681: dataIn1 = 32'd4
; 
32'd11682: dataIn1 = 32'd8
; 
32'd11683: dataIn1 = 32'd15
; 
32'd11684: dataIn1 = 32'd17
; 
32'd11685: dataIn1 = 32'd38
; 
32'd11686: dataIn1 = 32'd47
; 
32'd11687: dataIn1 = 32'd53
; 
32'd11688: dataIn1 = 32'd62
; 
32'd11689: dataIn1 = 32'd6
; 
32'd11690: dataIn1 = 32'd19
; 
32'd11691: dataIn1 = 32'd20
; 
32'd11692: dataIn1 = 32'd28
; 
32'd11693: dataIn1 = 32'd31
; 
32'd11694: dataIn1 = 32'd41
; 
32'd11695: dataIn1 = 32'd61
; 
32'd11696: dataIn1 = 32'd63
; 
32'd11697: dataIn1 = 32'd3
; 
32'd11698: dataIn1 = 32'd9
; 
32'd11699: dataIn1 = 32'd10
; 
32'd11700: dataIn1 = 32'd16
; 
32'd11701: dataIn1 = 32'd19
; 
32'd11702: dataIn1 = 32'd24
; 
32'd11703: dataIn1 = 32'd26
; 
32'd11704: dataIn1 = 32'd31
; 
32'd11705: dataIn1 = 32'd34
; 
32'd11706: dataIn1 = 32'd40
; 
32'd11707: dataIn1 = 32'd43
; 
32'd11708: dataIn1 = 32'd52
; 
32'd11709: dataIn1 = 32'd58
; 
32'd11710: dataIn1 = 32'd1
; 
32'd11711: dataIn1 = 32'd3
; 
32'd11712: dataIn1 = 32'd7
; 
32'd11713: dataIn1 = 32'd10
; 
32'd11714: dataIn1 = 32'd13
; 
32'd11715: dataIn1 = 32'd21
; 
32'd11716: dataIn1 = 32'd28
; 
32'd11717: dataIn1 = 32'd34
; 
32'd11718: dataIn1 = 32'd36
; 
32'd11719: dataIn1 = 32'd41
; 
32'd11720: dataIn1 = 32'd49
; 
32'd11721: dataIn1 = 32'd56
; 
32'd11722: dataIn1 = 32'd57
; 
32'd11723: dataIn1 = 32'd58
; 
32'd11724: dataIn1 = 32'd4
; 
32'd11725: dataIn1 = 32'd16
; 
32'd11726: dataIn1 = 32'd29
; 
32'd11727: dataIn1 = 32'd31
; 
32'd11728: dataIn1 = 32'd39
; 
32'd11729: dataIn1 = 32'd42
; 
32'd11730: dataIn1 = 32'd43
; 
32'd11731: dataIn1 = 32'd46
; 
32'd11732: dataIn1 = 32'd52
; 
32'd11733: dataIn1 = 32'd3
; 
32'd11734: dataIn1 = 32'd4
; 
32'd11735: dataIn1 = 32'd6
; 
32'd11736: dataIn1 = 32'd8
; 
32'd11737: dataIn1 = 32'd13
; 
32'd11738: dataIn1 = 32'd15
; 
32'd11739: dataIn1 = 32'd22
; 
32'd11740: dataIn1 = 32'd29
; 
32'd11741: dataIn1 = 32'd31
; 
32'd11742: dataIn1 = 32'd34
; 
32'd11743: dataIn1 = 32'd35
; 
32'd11744: dataIn1 = 32'd50
; 
32'd11745: dataIn1 = 32'd56
; 
32'd11746: dataIn1 = 32'd57
; 
32'd11747: dataIn1 = 32'd61
; 
32'd11748: dataIn1 = 32'd63
; 
32'd11749: dataIn1 = 32'd2
; 
32'd11750: dataIn1 = 32'd5
; 
32'd11751: dataIn1 = 32'd7
; 
32'd11752: dataIn1 = 32'd12
; 
32'd11753: dataIn1 = 32'd14
; 
32'd11754: dataIn1 = 32'd23
; 
32'd11755: dataIn1 = 32'd24
; 
32'd11756: dataIn1 = 32'd29
; 
32'd11757: dataIn1 = 32'd32
; 
32'd11758: dataIn1 = 32'd35
; 
32'd11759: dataIn1 = 32'd36
; 
32'd11760: dataIn1 = 32'd37
; 
32'd11761: dataIn1 = 32'd40
; 
32'd11762: dataIn1 = 32'd44
; 
32'd11763: dataIn1 = 32'd45
; 
32'd11764: dataIn1 = 32'd51
; 
32'd11765: dataIn1 = 32'd54
; 
32'd11766: dataIn1 = 32'd57
; 
32'd11767: dataIn1 = 32'd7
; 
32'd11768: dataIn1 = 32'd22
; 
32'd11769: dataIn1 = 32'd23
; 
32'd11770: dataIn1 = 32'd27
; 
32'd11771: dataIn1 = 32'd33
; 
32'd11772: dataIn1 = 32'd52
; 
32'd11773: dataIn1 = 32'd54
; 
32'd11774: dataIn1 = 32'd55
; 
32'd11775: dataIn1 = 32'd58
; 
32'd11776: dataIn1 = 32'd0
; 
32'd11777: dataIn1 = 32'd13
; 
32'd11778: dataIn1 = 32'd23
; 
32'd11779: dataIn1 = 32'd24
; 
32'd11780: dataIn1 = 32'd25
; 
32'd11781: dataIn1 = 32'd27
; 
32'd11782: dataIn1 = 32'd33
; 
32'd11783: dataIn1 = 32'd42
; 
32'd11784: dataIn1 = 32'd44
; 
32'd11785: dataIn1 = 32'd50
; 
32'd11786: dataIn1 = 32'd51
; 
32'd11787: dataIn1 = 32'd54
; 
32'd11788: dataIn1 = 32'd56
; 
32'd11789: dataIn1 = 32'd57
; 
32'd11790: dataIn1 = 32'd60
; 
32'd11791: dataIn1 = 32'd4
; 
32'd11792: dataIn1 = 32'd17
; 
32'd11793: dataIn1 = 32'd19
; 
32'd11794: dataIn1 = 32'd28
; 
32'd11795: dataIn1 = 32'd34
; 
32'd11796: dataIn1 = 32'd38
; 
32'd11797: dataIn1 = 32'd42
; 
32'd11798: dataIn1 = 32'd46
; 
32'd11799: dataIn1 = 32'd48
; 
32'd11800: dataIn1 = 32'd57
; 
32'd11801: dataIn1 = 32'd3
; 
32'd11802: dataIn1 = 32'd4
; 
32'd11803: dataIn1 = 32'd6
; 
32'd11804: dataIn1 = 32'd7
; 
32'd11805: dataIn1 = 32'd14
; 
32'd11806: dataIn1 = 32'd18
; 
32'd11807: dataIn1 = 32'd19
; 
32'd11808: dataIn1 = 32'd22
; 
32'd11809: dataIn1 = 32'd34
; 
32'd11810: dataIn1 = 32'd46
; 
32'd11811: dataIn1 = 32'd60
; 
32'd11812: dataIn1 = 32'd1
; 
32'd11813: dataIn1 = 32'd5
; 
32'd11814: dataIn1 = 32'd6
; 
32'd11815: dataIn1 = 32'd7
; 
32'd11816: dataIn1 = 32'd11
; 
32'd11817: dataIn1 = 32'd21
; 
32'd11818: dataIn1 = 32'd26
; 
32'd11819: dataIn1 = 32'd28
; 
32'd11820: dataIn1 = 32'd32
; 
32'd11821: dataIn1 = 32'd33
; 
32'd11822: dataIn1 = 32'd36
; 
32'd11823: dataIn1 = 32'd38
; 
32'd11824: dataIn1 = 32'd41
; 
32'd11825: dataIn1 = 32'd45
; 
32'd11826: dataIn1 = 32'd1
; 
32'd11827: dataIn1 = 32'd3
; 
32'd11828: dataIn1 = 32'd9
; 
32'd11829: dataIn1 = 32'd10
; 
32'd11830: dataIn1 = 32'd13
; 
32'd11831: dataIn1 = 32'd18
; 
32'd11832: dataIn1 = 32'd29
; 
32'd11833: dataIn1 = 32'd30
; 
32'd11834: dataIn1 = 32'd35
; 
32'd11835: dataIn1 = 32'd39
; 
32'd11836: dataIn1 = 32'd42
; 
32'd11837: dataIn1 = 32'd46
; 
32'd11838: dataIn1 = 32'd49
; 
32'd11839: dataIn1 = 32'd50
; 
32'd11840: dataIn1 = 32'd51
; 
32'd11841: dataIn1 = 32'd52
; 
32'd11842: dataIn1 = 32'd1
; 
32'd11843: dataIn1 = 32'd12
; 
32'd11844: dataIn1 = 32'd13
; 
32'd11845: dataIn1 = 32'd17
; 
32'd11846: dataIn1 = 32'd21
; 
32'd11847: dataIn1 = 32'd24
; 
32'd11848: dataIn1 = 32'd34
; 
32'd11849: dataIn1 = 32'd38
; 
32'd11850: dataIn1 = 32'd39
; 
32'd11851: dataIn1 = 32'd40
; 
32'd11852: dataIn1 = 32'd42
; 
32'd11853: dataIn1 = 32'd45
; 
32'd11854: dataIn1 = 32'd46
; 
32'd11855: dataIn1 = 32'd47
; 
32'd11856: dataIn1 = 32'd53
; 
32'd11857: dataIn1 = 32'd0
; 
32'd11858: dataIn1 = 32'd4
; 
32'd11859: dataIn1 = 32'd9
; 
32'd11860: dataIn1 = 32'd12
; 
32'd11861: dataIn1 = 32'd14
; 
32'd11862: dataIn1 = 32'd25
; 
32'd11863: dataIn1 = 32'd27
; 
32'd11864: dataIn1 = 32'd30
; 
32'd11865: dataIn1 = 32'd31
; 
32'd11866: dataIn1 = 32'd35
; 
32'd11867: dataIn1 = 32'd36
; 
32'd11868: dataIn1 = 32'd53
; 
32'd11869: dataIn1 = 32'd56
; 
32'd11870: dataIn1 = 32'd59
; 
32'd11871: dataIn1 = 32'd61
; 
32'd11872: dataIn1 = 32'd13
; 
32'd11873: dataIn1 = 32'd14
; 
32'd11874: dataIn1 = 32'd15
; 
32'd11875: dataIn1 = 32'd22
; 
32'd11876: dataIn1 = 32'd23
; 
32'd11877: dataIn1 = 32'd28
; 
32'd11878: dataIn1 = 32'd35
; 
32'd11879: dataIn1 = 32'd36
; 
32'd11880: dataIn1 = 32'd43
; 
32'd11881: dataIn1 = 32'd44
; 
32'd11882: dataIn1 = 32'd46
; 
32'd11883: dataIn1 = 32'd50
; 
32'd11884: dataIn1 = 32'd52
; 
32'd11885: dataIn1 = 32'd55
; 
32'd11886: dataIn1 = 32'd62
; 
32'd11887: dataIn1 = 32'd63
; 
32'd11888: dataIn1 = 32'd2
; 
32'd11889: dataIn1 = 32'd4
; 
32'd11890: dataIn1 = 32'd5
; 
32'd11891: dataIn1 = 32'd8
; 
32'd11892: dataIn1 = 32'd11
; 
32'd11893: dataIn1 = 32'd16
; 
32'd11894: dataIn1 = 32'd19
; 
32'd11895: dataIn1 = 32'd23
; 
32'd11896: dataIn1 = 32'd29
; 
32'd11897: dataIn1 = 32'd31
; 
32'd11898: dataIn1 = 32'd32
; 
32'd11899: dataIn1 = 32'd33
; 
32'd11900: dataIn1 = 32'd45
; 
32'd11901: dataIn1 = 32'd50
; 
32'd11902: dataIn1 = 32'd51
; 
32'd11903: dataIn1 = 32'd58
; 
32'd11904: dataIn1 = 32'd61
; 
32'd11905: dataIn1 = 32'd63
; 
32'd11906: dataIn1 = 32'd6
; 
32'd11907: dataIn1 = 32'd12
; 
32'd11908: dataIn1 = 32'd18
; 
32'd11909: dataIn1 = 32'd24
; 
32'd11910: dataIn1 = 32'd33
; 
32'd11911: dataIn1 = 32'd34
; 
32'd11912: dataIn1 = 32'd41
; 
32'd11913: dataIn1 = 32'd42
; 
32'd11914: dataIn1 = 32'd59
; 
32'd11915: dataIn1 = 32'd60
; 
32'd11916: dataIn1 = 32'd14
; 
32'd11917: dataIn1 = 32'd21
; 
32'd11918: dataIn1 = 32'd22
; 
32'd11919: dataIn1 = 32'd25
; 
32'd11920: dataIn1 = 32'd27
; 
32'd11921: dataIn1 = 32'd28
; 
32'd11922: dataIn1 = 32'd38
; 
32'd11923: dataIn1 = 32'd60
; 
32'd11924: dataIn1 = 32'd62
; 
32'd11925: dataIn1 = 32'd4
; 
32'd11926: dataIn1 = 32'd7
; 
32'd11927: dataIn1 = 32'd17
; 
32'd11928: dataIn1 = 32'd31
; 
32'd11929: dataIn1 = 32'd39
; 
32'd11930: dataIn1 = 32'd43
; 
32'd11931: dataIn1 = 32'd50
; 
32'd11932: dataIn1 = 32'd51
; 
32'd11933: dataIn1 = 32'd57
; 
32'd11934: dataIn1 = 32'd61
; 
32'd11935: dataIn1 = 32'd1
; 
32'd11936: dataIn1 = 32'd3
; 
32'd11937: dataIn1 = 32'd10
; 
32'd11938: dataIn1 = 32'd17
; 
32'd11939: dataIn1 = 32'd26
; 
32'd11940: dataIn1 = 32'd31
; 
32'd11941: dataIn1 = 32'd33
; 
32'd11942: dataIn1 = 32'd42
; 
32'd11943: dataIn1 = 32'd49
; 
32'd11944: dataIn1 = 32'd55
; 
32'd11945: dataIn1 = 32'd58
; 
32'd11946: dataIn1 = 32'd0
; 
32'd11947: dataIn1 = 32'd13
; 
32'd11948: dataIn1 = 32'd15
; 
32'd11949: dataIn1 = 32'd32
; 
32'd11950: dataIn1 = 32'd42
; 
32'd11951: dataIn1 = 32'd51
; 
32'd11952: dataIn1 = 32'd54
; 
32'd11953: dataIn1 = 32'd55
; 
32'd11954: dataIn1 = 32'd59
; 
32'd11955: dataIn1 = 32'd5
; 
32'd11956: dataIn1 = 32'd9
; 
32'd11957: dataIn1 = 32'd25
; 
32'd11958: dataIn1 = 32'd30
; 
32'd11959: dataIn1 = 32'd34
; 
32'd11960: dataIn1 = 32'd37
; 
32'd11961: dataIn1 = 32'd40
; 
32'd11962: dataIn1 = 32'd47
; 
32'd11963: dataIn1 = 32'd48
; 
32'd11964: dataIn1 = 32'd55
; 
32'd11965: dataIn1 = 32'd56
; 
32'd11966: dataIn1 = 32'd60
; 
32'd11967: dataIn1 = 32'd63
; 
32'd11968: dataIn1 = 32'd0
; 
32'd11969: dataIn1 = 32'd1
; 
32'd11970: dataIn1 = 32'd4
; 
32'd11971: dataIn1 = 32'd6
; 
32'd11972: dataIn1 = 32'd9
; 
32'd11973: dataIn1 = 32'd10
; 
32'd11974: dataIn1 = 32'd19
; 
32'd11975: dataIn1 = 32'd20
; 
32'd11976: dataIn1 = 32'd21
; 
32'd11977: dataIn1 = 32'd28
; 
32'd11978: dataIn1 = 32'd31
; 
32'd11979: dataIn1 = 32'd37
; 
32'd11980: dataIn1 = 32'd40
; 
32'd11981: dataIn1 = 32'd42
; 
32'd11982: dataIn1 = 32'd47
; 
32'd11983: dataIn1 = 32'd49
; 
32'd11984: dataIn1 = 32'd53
; 
32'd11985: dataIn1 = 32'd54
; 
32'd11986: dataIn1 = 32'd57
; 
32'd11987: dataIn1 = 32'd2
; 
32'd11988: dataIn1 = 32'd8
; 
32'd11989: dataIn1 = 32'd20
; 
32'd11990: dataIn1 = 32'd26
; 
32'd11991: dataIn1 = 32'd29
; 
32'd11992: dataIn1 = 32'd32
; 
32'd11993: dataIn1 = 32'd37
; 
32'd11994: dataIn1 = 32'd38
; 
32'd11995: dataIn1 = 32'd44
; 
32'd11996: dataIn1 = 32'd48
; 
32'd11997: dataIn1 = 32'd49
; 
32'd11998: dataIn1 = 32'd57
; 
32'd11999: dataIn1 = 32'd62
; 
32'd12000: dataIn1 = 32'd1
; 
32'd12001: dataIn1 = 32'd3
; 
32'd12002: dataIn1 = 32'd15
; 
32'd12003: dataIn1 = 32'd20
; 
32'd12004: dataIn1 = 32'd31
; 
32'd12005: dataIn1 = 32'd33
; 
32'd12006: dataIn1 = 32'd37
; 
32'd12007: dataIn1 = 32'd41
; 
32'd12008: dataIn1 = 32'd48
; 
32'd12009: dataIn1 = 32'd53
; 
32'd12010: dataIn1 = 32'd54
; 
32'd12011: dataIn1 = 32'd58
; 
32'd12012: dataIn1 = 32'd62
; 
32'd12013: dataIn1 = 32'd2
; 
32'd12014: dataIn1 = 32'd14
; 
32'd12015: dataIn1 = 32'd19
; 
32'd12016: dataIn1 = 32'd21
; 
32'd12017: dataIn1 = 32'd31
; 
32'd12018: dataIn1 = 32'd42
; 
32'd12019: dataIn1 = 32'd44
; 
32'd12020: dataIn1 = 32'd45
; 
32'd12021: dataIn1 = 32'd46
; 
32'd12022: dataIn1 = 32'd51
; 
32'd12023: dataIn1 = 32'd52
; 
32'd12024: dataIn1 = 32'd55
; 
32'd12025: dataIn1 = 32'd57
; 
32'd12026: dataIn1 = 32'd60
; 
32'd12027: dataIn1 = 32'd12
; 
32'd12028: dataIn1 = 32'd19
; 
32'd12029: dataIn1 = 32'd20
; 
32'd12030: dataIn1 = 32'd22
; 
32'd12031: dataIn1 = 32'd35
; 
32'd12032: dataIn1 = 32'd36
; 
32'd12033: dataIn1 = 32'd41
; 
32'd12034: dataIn1 = 32'd49
; 
32'd12035: dataIn1 = 32'd53
; 
32'd12036: dataIn1 = 32'd59
; 
32'd12037: dataIn1 = 32'd60
; 
32'd12038: dataIn1 = 32'd3
; 
32'd12039: dataIn1 = 32'd20
; 
32'd12040: dataIn1 = 32'd22
; 
32'd12041: dataIn1 = 32'd25
; 
32'd12042: dataIn1 = 32'd26
; 
32'd12043: dataIn1 = 32'd31
; 
32'd12044: dataIn1 = 32'd35
; 
32'd12045: dataIn1 = 32'd38
; 
32'd12046: dataIn1 = 32'd42
; 
32'd12047: dataIn1 = 32'd45
; 
32'd12048: dataIn1 = 32'd48
; 
32'd12049: dataIn1 = 32'd53
; 
32'd12050: dataIn1 = 32'd1
; 
32'd12051: dataIn1 = 32'd3
; 
32'd12052: dataIn1 = 32'd10
; 
32'd12053: dataIn1 = 32'd11
; 
32'd12054: dataIn1 = 32'd25
; 
32'd12055: dataIn1 = 32'd39
; 
32'd12056: dataIn1 = 32'd42
; 
32'd12057: dataIn1 = 32'd43
; 
32'd12058: dataIn1 = 32'd52
; 
32'd12059: dataIn1 = 32'd3
; 
32'd12060: dataIn1 = 32'd4
; 
32'd12061: dataIn1 = 32'd5
; 
32'd12062: dataIn1 = 32'd9
; 
32'd12063: dataIn1 = 32'd10
; 
32'd12064: dataIn1 = 32'd14
; 
32'd12065: dataIn1 = 32'd18
; 
32'd12066: dataIn1 = 32'd19
; 
32'd12067: dataIn1 = 32'd23
; 
32'd12068: dataIn1 = 32'd26
; 
32'd12069: dataIn1 = 32'd31
; 
32'd12070: dataIn1 = 32'd38
; 
32'd12071: dataIn1 = 32'd42
; 
32'd12072: dataIn1 = 32'd47
; 
32'd12073: dataIn1 = 32'd56
; 
32'd12074: dataIn1 = 32'd57
; 
32'd12075: dataIn1 = 32'd60
; 
32'd12076: dataIn1 = 32'd4
; 
32'd12077: dataIn1 = 32'd7
; 
32'd12078: dataIn1 = 32'd12
; 
32'd12079: dataIn1 = 32'd14
; 
32'd12080: dataIn1 = 32'd25
; 
32'd12081: dataIn1 = 32'd26
; 
32'd12082: dataIn1 = 32'd40
; 
32'd12083: dataIn1 = 32'd45
; 
32'd12084: dataIn1 = 32'd52
; 
32'd12085: dataIn1 = 32'd57
; 
32'd12086: dataIn1 = 32'd61
; 
32'd12087: dataIn1 = 32'd62
; 
32'd12088: dataIn1 = 32'd6
; 
32'd12089: dataIn1 = 32'd12
; 
32'd12090: dataIn1 = 32'd17
; 
32'd12091: dataIn1 = 32'd25
; 
32'd12092: dataIn1 = 32'd37
; 
32'd12093: dataIn1 = 32'd38
; 
32'd12094: dataIn1 = 32'd40
; 
32'd12095: dataIn1 = 32'd43
; 
32'd12096: dataIn1 = 32'd44
; 
32'd12097: dataIn1 = 32'd61
; 
32'd12098: dataIn1 = 32'd63
; 
32'd12099: dataIn1 = 32'd7
; 
32'd12100: dataIn1 = 32'd14
; 
32'd12101: dataIn1 = 32'd22
; 
32'd12102: dataIn1 = 32'd24
; 
32'd12103: dataIn1 = 32'd41
; 
32'd12104: dataIn1 = 32'd44
; 
32'd12105: dataIn1 = 32'd45
; 
32'd12106: dataIn1 = 32'd58
; 
32'd12107: dataIn1 = 32'd61
; 
32'd12108: dataIn1 = 32'd3
; 
32'd12109: dataIn1 = 32'd11
; 
32'd12110: dataIn1 = 32'd13
; 
32'd12111: dataIn1 = 32'd22
; 
32'd12112: dataIn1 = 32'd25
; 
32'd12113: dataIn1 = 32'd30
; 
32'd12114: dataIn1 = 32'd31
; 
32'd12115: dataIn1 = 32'd40
; 
32'd12116: dataIn1 = 32'd41
; 
32'd12117: dataIn1 = 32'd43
; 
32'd12118: dataIn1 = 32'd46
; 
32'd12119: dataIn1 = 32'd53
; 
32'd12120: dataIn1 = 32'd58
; 
32'd12121: dataIn1 = 32'd2
; 
32'd12122: dataIn1 = 32'd3
; 
32'd12123: dataIn1 = 32'd9
; 
32'd12124: dataIn1 = 32'd14
; 
32'd12125: dataIn1 = 32'd15
; 
32'd12126: dataIn1 = 32'd17
; 
32'd12127: dataIn1 = 32'd18
; 
32'd12128: dataIn1 = 32'd20
; 
32'd12129: dataIn1 = 32'd27
; 
32'd12130: dataIn1 = 32'd29
; 
32'd12131: dataIn1 = 32'd31
; 
32'd12132: dataIn1 = 32'd32
; 
32'd12133: dataIn1 = 32'd37
; 
32'd12134: dataIn1 = 32'd43
; 
32'd12135: dataIn1 = 32'd4
; 
32'd12136: dataIn1 = 32'd5
; 
32'd12137: dataIn1 = 32'd11
; 
32'd12138: dataIn1 = 32'd13
; 
32'd12139: dataIn1 = 32'd30
; 
32'd12140: dataIn1 = 32'd34
; 
32'd12141: dataIn1 = 32'd35
; 
32'd12142: dataIn1 = 32'd36
; 
32'd12143: dataIn1 = 32'd43
; 
32'd12144: dataIn1 = 32'd46
; 
32'd12145: dataIn1 = 32'd57
; 
32'd12146: dataIn1 = 32'd61
; 
32'd12147: dataIn1 = 32'd63
; 
32'd12148: dataIn1 = 32'd0
; 
32'd12149: dataIn1 = 32'd1
; 
32'd12150: dataIn1 = 32'd3
; 
32'd12151: dataIn1 = 32'd9
; 
32'd12152: dataIn1 = 32'd17
; 
32'd12153: dataIn1 = 32'd21
; 
32'd12154: dataIn1 = 32'd24
; 
32'd12155: dataIn1 = 32'd26
; 
32'd12156: dataIn1 = 32'd33
; 
32'd12157: dataIn1 = 32'd39
; 
32'd12158: dataIn1 = 32'd42
; 
32'd12159: dataIn1 = 32'd50
; 
32'd12160: dataIn1 = 32'd59
; 
32'd12161: dataIn1 = 32'd63
; 
32'd12162: dataIn1 = 32'd4
; 
32'd12163: dataIn1 = 32'd7
; 
32'd12164: dataIn1 = 32'd28
; 
32'd12165: dataIn1 = 32'd29
; 
32'd12166: dataIn1 = 32'd36
; 
32'd12167: dataIn1 = 32'd38
; 
32'd12168: dataIn1 = 32'd40
; 
32'd12169: dataIn1 = 32'd41
; 
32'd12170: dataIn1 = 32'd55
; 
32'd12171: dataIn1 = 32'd3
; 
32'd12172: dataIn1 = 32'd4
; 
32'd12173: dataIn1 = 32'd14
; 
32'd12174: dataIn1 = 32'd16
; 
32'd12175: dataIn1 = 32'd23
; 
32'd12176: dataIn1 = 32'd31
; 
32'd12177: dataIn1 = 32'd34
; 
32'd12178: dataIn1 = 32'd44
; 
32'd12179: dataIn1 = 32'd54
; 
32'd12180: dataIn1 = 32'd63
; 
32'd12181: dataIn1 = 32'd0
; 
32'd12182: dataIn1 = 32'd3
; 
32'd12183: dataIn1 = 32'd4
; 
32'd12184: dataIn1 = 32'd5
; 
32'd12185: dataIn1 = 32'd6
; 
32'd12186: dataIn1 = 32'd8
; 
32'd12187: dataIn1 = 32'd9
; 
32'd12188: dataIn1 = 32'd12
; 
32'd12189: dataIn1 = 32'd20
; 
32'd12190: dataIn1 = 32'd26
; 
32'd12191: dataIn1 = 32'd43
; 
32'd12192: dataIn1 = 32'd45
; 
32'd12193: dataIn1 = 32'd46
; 
32'd12194: dataIn1 = 32'd1
; 
32'd12195: dataIn1 = 32'd12
; 
32'd12196: dataIn1 = 32'd17
; 
32'd12197: dataIn1 = 32'd27
; 
32'd12198: dataIn1 = 32'd32
; 
32'd12199: dataIn1 = 32'd36
; 
32'd12200: dataIn1 = 32'd38
; 
32'd12201: dataIn1 = 32'd41
; 
32'd12202: dataIn1 = 32'd42
; 
32'd12203: dataIn1 = 32'd53
; 
32'd12204: dataIn1 = 32'd54
; 
32'd12205: dataIn1 = 32'd55
; 
32'd12206: dataIn1 = 32'd61
; 
32'd12207: dataIn1 = 32'd0
; 
32'd12208: dataIn1 = 32'd1
; 
32'd12209: dataIn1 = 32'd2
; 
32'd12210: dataIn1 = 32'd3
; 
32'd12211: dataIn1 = 32'd14
; 
32'd12212: dataIn1 = 32'd15
; 
32'd12213: dataIn1 = 32'd22
; 
32'd12214: dataIn1 = 32'd24
; 
32'd12215: dataIn1 = 32'd30
; 
32'd12216: dataIn1 = 32'd32
; 
32'd12217: dataIn1 = 32'd34
; 
32'd12218: dataIn1 = 32'd38
; 
32'd12219: dataIn1 = 32'd41
; 
32'd12220: dataIn1 = 32'd42
; 
32'd12221: dataIn1 = 32'd44
; 
32'd12222: dataIn1 = 32'd47
; 
32'd12223: dataIn1 = 32'd58
; 
32'd12224: dataIn1 = 32'd59
; 
32'd12225: dataIn1 = 32'd62
; 
32'd12226: dataIn1 = 32'd0
; 
32'd12227: dataIn1 = 32'd1
; 
32'd12228: dataIn1 = 32'd4
; 
32'd12229: dataIn1 = 32'd5
; 
32'd12230: dataIn1 = 32'd15
; 
32'd12231: dataIn1 = 32'd17
; 
32'd12232: dataIn1 = 32'd20
; 
32'd12233: dataIn1 = 32'd31
; 
32'd12234: dataIn1 = 32'd34
; 
32'd12235: dataIn1 = 32'd36
; 
32'd12236: dataIn1 = 32'd40
; 
32'd12237: dataIn1 = 32'd41
; 
32'd12238: dataIn1 = 32'd59
; 
32'd12239: dataIn1 = 32'd60
; 
32'd12240: dataIn1 = 32'd61
; 
32'd12241: dataIn1 = 32'd63
; 
32'd12242: dataIn1 = 32'd0
; 
32'd12243: dataIn1 = 32'd2
; 
32'd12244: dataIn1 = 32'd3
; 
32'd12245: dataIn1 = 32'd10
; 
32'd12246: dataIn1 = 32'd14
; 
32'd12247: dataIn1 = 32'd17
; 
32'd12248: dataIn1 = 32'd19
; 
32'd12249: dataIn1 = 32'd25
; 
32'd12250: dataIn1 = 32'd42
; 
32'd12251: dataIn1 = 32'd53
; 
32'd12252: dataIn1 = 32'd58
; 
32'd12253: dataIn1 = 32'd60
; 
32'd12254: dataIn1 = 32'd1
; 
32'd12255: dataIn1 = 32'd5
; 
32'd12256: dataIn1 = 32'd7
; 
32'd12257: dataIn1 = 32'd15
; 
32'd12258: dataIn1 = 32'd17
; 
32'd12259: dataIn1 = 32'd24
; 
32'd12260: dataIn1 = 32'd25
; 
32'd12261: dataIn1 = 32'd26
; 
32'd12262: dataIn1 = 32'd33
; 
32'd12263: dataIn1 = 32'd50
; 
32'd12264: dataIn1 = 32'd53
; 
32'd12265: dataIn1 = 32'd3
; 
32'd12266: dataIn1 = 32'd15
; 
32'd12267: dataIn1 = 32'd18
; 
32'd12268: dataIn1 = 32'd23
; 
32'd12269: dataIn1 = 32'd27
; 
32'd12270: dataIn1 = 32'd28
; 
32'd12271: dataIn1 = 32'd36
; 
32'd12272: dataIn1 = 32'd38
; 
32'd12273: dataIn1 = 32'd47
; 
32'd12274: dataIn1 = 32'd48
; 
32'd12275: dataIn1 = 32'd51
; 
32'd12276: dataIn1 = 32'd8
; 
32'd12277: dataIn1 = 32'd10
; 
32'd12278: dataIn1 = 32'd13
; 
32'd12279: dataIn1 = 32'd14
; 
32'd12280: dataIn1 = 32'd15
; 
32'd12281: dataIn1 = 32'd24
; 
32'd12282: dataIn1 = 32'd25
; 
32'd12283: dataIn1 = 32'd30
; 
32'd12284: dataIn1 = 32'd37
; 
32'd12285: dataIn1 = 32'd47
; 
32'd12286: dataIn1 = 32'd53
; 
32'd12287: dataIn1 = 32'd56
; 
32'd12288: dataIn1 = 32'd59
; 
32'd12289: dataIn1 = 32'd0
; 
32'd12290: dataIn1 = 32'd16
; 
32'd12291: dataIn1 = 32'd18
; 
32'd12292: dataIn1 = 32'd25
; 
32'd12293: dataIn1 = 32'd27
; 
32'd12294: dataIn1 = 32'd35
; 
32'd12295: dataIn1 = 32'd37
; 
32'd12296: dataIn1 = 32'd40
; 
32'd12297: dataIn1 = 32'd42
; 
32'd12298: dataIn1 = 32'd44
; 
32'd12299: dataIn1 = 32'd50
; 
32'd12300: dataIn1 = 32'd58
; 
32'd12301: dataIn1 = 32'd60
; 
32'd12302: dataIn1 = 32'd8
; 
32'd12303: dataIn1 = 32'd20
; 
32'd12304: dataIn1 = 32'd21
; 
32'd12305: dataIn1 = 32'd33
; 
32'd12306: dataIn1 = 32'd37
; 
32'd12307: dataIn1 = 32'd38
; 
32'd12308: dataIn1 = 32'd48
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd88; 
32'd3: dataIn2 = 32'd36; 
32'd4: dataIn2 = 32'd16; 
32'd5: dataIn2 = 32'd42; 
32'd6: dataIn2 = 32'd2; 
32'd7: dataIn2 = 32'd47; 
32'd8: dataIn2 = 32'd57; 
32'd9: dataIn2 = 32'd10; 
32'd10: dataIn2 = 32'd12; 
32'd11: dataIn2 = 32'd46; 
32'd12: dataIn2 = 32'd47; 
32'd13: dataIn2 = 32'd29; 
32'd14: dataIn2 = 32'd74; 
32'd15: dataIn2 = 32'd7; 
32'd16: dataIn2 = 32'd63; 
32'd17: dataIn2 = 32'd23; 
32'd18: dataIn2 = 32'd14; 
32'd19: dataIn2 = 32'd37; 
32'd20: dataIn2 = 32'd51; 
32'd21: dataIn2 = 32'd48; 
32'd22: dataIn2 = 32'd95; 
32'd23: dataIn2 = 32'd87; 
32'd24: dataIn2 = 32'd78; 
32'd25: dataIn2 = 32'd5; 
32'd26: dataIn2 = 32'd66; 
32'd27: dataIn2 = 32'd71; 
32'd28: dataIn2 = 32'd75; 
32'd29: dataIn2 = 32'd25; 
32'd30: dataIn2 = 32'd74; 
32'd31: dataIn2 = 32'd78; 
32'd32: dataIn2 = 32'd31; 
32'd33: dataIn2 = 32'd39; 
32'd34: dataIn2 = 32'd28; 
32'd35: dataIn2 = 32'd23; 
32'd36: dataIn2 = 32'd83; 
32'd37: dataIn2 = 32'd55; 
32'd38: dataIn2 = 32'd55; 
32'd39: dataIn2 = 32'd100; 
32'd40: dataIn2 = 32'd22; 
32'd41: dataIn2 = 32'd47; 
32'd42: dataIn2 = 32'd9; 
32'd43: dataIn2 = 32'd90; 
32'd44: dataIn2 = 32'd63; 
32'd45: dataIn2 = 32'd45; 
32'd46: dataIn2 = 32'd14; 
32'd47: dataIn2 = 32'd49; 
32'd48: dataIn2 = 32'd37; 
32'd49: dataIn2 = 32'd93; 
32'd50: dataIn2 = 32'd6; 
32'd51: dataIn2 = 32'd1; 
32'd52: dataIn2 = 32'd4; 
32'd53: dataIn2 = 32'd30; 
32'd54: dataIn2 = 32'd89; 
32'd55: dataIn2 = 32'd47; 
32'd56: dataIn2 = 32'd61; 
32'd57: dataIn2 = 32'd74; 
32'd58: dataIn2 = 32'd40; 
32'd59: dataIn2 = 32'd27; 
32'd60: dataIn2 = 32'd72; 
32'd61: dataIn2 = 32'd49; 
32'd62: dataIn2 = 32'd77; 
32'd63: dataIn2 = 32'd36; 
32'd64: dataIn2 = 32'd89; 
32'd65: dataIn2 = 32'd32; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd330: dataIn2 = 32'd92; 
32'd331: dataIn2 = 32'd50; 
32'd332: dataIn2 = 32'd36; 
32'd333: dataIn2 = 32'd67; 
32'd334: dataIn2 = 32'd95; 
32'd335: dataIn2 = 32'd96; 
32'd336: dataIn2 = 32'd77; 
32'd337: dataIn2 = 32'd80; 
32'd338: dataIn2 = 32'd27; 
32'd339: dataIn2 = 32'd65; 
32'd340: dataIn2 = 32'd84; 
32'd341: dataIn2 = 32'd30; 
32'd342: dataIn2 = 32'd92; 
32'd343: dataIn2 = 32'd96; 
32'd344: dataIn2 = 32'd93; 
32'd345: dataIn2 = 32'd81; 
32'd346: dataIn2 = 32'd89; 
32'd347: dataIn2 = 32'd18; 
32'd348: dataIn2 = 32'd59; 
32'd349: dataIn2 = 32'd60; 
32'd350: dataIn2 = 32'd30; 
32'd351: dataIn2 = 32'd55; 
32'd352: dataIn2 = 32'd78; 
32'd353: dataIn2 = 32'd61; 
32'd354: dataIn2 = 32'd89; 
32'd355: dataIn2 = 32'd75; 
32'd356: dataIn2 = 32'd42; 
32'd357: dataIn2 = 32'd79; 
32'd358: dataIn2 = 32'd23; 
32'd359: dataIn2 = 32'd73; 
32'd360: dataIn2 = 32'd45; 
32'd361: dataIn2 = 32'd78; 
32'd362: dataIn2 = 32'd63; 
32'd363: dataIn2 = 32'd75; 
32'd364: dataIn2 = 32'd41; 
32'd365: dataIn2 = 32'd71; 
32'd366: dataIn2 = 32'd52; 
32'd367: dataIn2 = 32'd61; 
32'd368: dataIn2 = 32'd53; 
32'd369: dataIn2 = 32'd69; 
32'd370: dataIn2 = 32'd21; 
32'd371: dataIn2 = 32'd10; 
32'd372: dataIn2 = 32'd11; 
32'd373: dataIn2 = 32'd44; 
32'd374: dataIn2 = 32'd28; 
32'd375: dataIn2 = 32'd4; 
32'd376: dataIn2 = 32'd35; 
32'd377: dataIn2 = 32'd49; 
32'd378: dataIn2 = 32'd69; 
32'd379: dataIn2 = 32'd83; 
32'd380: dataIn2 = 32'd38; 
32'd381: dataIn2 = 32'd79; 
32'd382: dataIn2 = 32'd35; 
32'd383: dataIn2 = 32'd87; 
32'd384: dataIn2 = 32'd68; 
32'd385: dataIn2 = 32'd91; 
32'd386: dataIn2 = 32'd60; 
32'd387: dataIn2 = 32'd100; 
32'd388: dataIn2 = 32'd100; 
32'd389: dataIn2 = 32'd54; 
32'd390: dataIn2 = 32'd28; 
32'd391: dataIn2 = 32'd70; 
32'd392: dataIn2 = 32'd70; 
32'd393: dataIn2 = 32'd30; 
32'd394: dataIn2 = 32'd77; 
32'd395: dataIn2 = 32'd74; 
32'd396: dataIn2 = 32'd69; 
32'd397: dataIn2 = 32'd56; 
32'd398: dataIn2 = 32'd48; 
32'd399: dataIn2 = 32'd28; 
32'd400: dataIn2 = 32'd93; 
32'd401: dataIn2 = 32'd33; 
32'd402: dataIn2 = 32'd4; 
32'd403: dataIn2 = 32'd53; 
32'd404: dataIn2 = 32'd58; 
32'd405: dataIn2 = 32'd79; 
32'd406: dataIn2 = 32'd83; 
32'd407: dataIn2 = 32'd88; 
32'd408: dataIn2 = 32'd56; 
32'd409: dataIn2 = 32'd28; 
32'd410: dataIn2 = 32'd76; 
32'd411: dataIn2 = 32'd0; 
32'd412: dataIn2 = 32'd31; 
32'd413: dataIn2 = 32'd10; 
32'd414: dataIn2 = 32'd100; 
32'd415: dataIn2 = 32'd51; 
32'd416: dataIn2 = 32'd61; 
32'd417: dataIn2 = 32'd37; 
32'd418: dataIn2 = 32'd81; 
32'd419: dataIn2 = 32'd71; 
32'd420: dataIn2 = 32'd19; 
32'd421: dataIn2 = 32'd97; 
32'd422: dataIn2 = 32'd70; 
32'd423: dataIn2 = 32'd55; 
32'd424: dataIn2 = 32'd87; 
32'd425: dataIn2 = 32'd86; 
32'd426: dataIn2 = 32'd97; 
32'd427: dataIn2 = 32'd79; 
32'd428: dataIn2 = 32'd18; 
32'd429: dataIn2 = 32'd80; 
32'd430: dataIn2 = 32'd87; 
32'd431: dataIn2 = 32'd28; 
32'd432: dataIn2 = 32'd41; 
32'd433: dataIn2 = 32'd88; 
32'd434: dataIn2 = 32'd86; 
32'd435: dataIn2 = 32'd58; 
32'd436: dataIn2 = 32'd19; 
32'd437: dataIn2 = 32'd52; 
32'd438: dataIn2 = 32'd98; 
32'd439: dataIn2 = 32'd85; 
32'd440: dataIn2 = 32'd42; 
32'd441: dataIn2 = 32'd74; 
32'd442: dataIn2 = 32'd38; 
32'd443: dataIn2 = 32'd41; 
32'd444: dataIn2 = 32'd0; 
32'd445: dataIn2 = 32'd15; 
32'd446: dataIn2 = 32'd89; 
32'd447: dataIn2 = 32'd47; 
32'd448: dataIn2 = 32'd81; 
32'd449: dataIn2 = 32'd84; 
32'd450: dataIn2 = 32'd37; 
32'd451: dataIn2 = 32'd88; 
32'd452: dataIn2 = 32'd56; 
32'd453: dataIn2 = 32'd13; 
32'd454: dataIn2 = 32'd87; 
32'd455: dataIn2 = 32'd64; 
32'd456: dataIn2 = 32'd41; 
32'd457: dataIn2 = 32'd69; 
32'd458: dataIn2 = 32'd52; 
32'd459: dataIn2 = 32'd98; 
32'd460: dataIn2 = 32'd88; 
32'd461: dataIn2 = 32'd67; 
32'd462: dataIn2 = 32'd26; 
32'd463: dataIn2 = 32'd11; 
32'd464: dataIn2 = 32'd25; 
32'd465: dataIn2 = 32'd18; 
32'd466: dataIn2 = 32'd2; 
32'd467: dataIn2 = 32'd20; 
32'd468: dataIn2 = 32'd27; 
32'd469: dataIn2 = 32'd99; 
32'd470: dataIn2 = 32'd45; 
32'd471: dataIn2 = 32'd55; 
32'd472: dataIn2 = 32'd45; 
32'd473: dataIn2 = 32'd57; 
32'd474: dataIn2 = 32'd42; 
32'd475: dataIn2 = 32'd95; 
32'd476: dataIn2 = 32'd19; 
32'd477: dataIn2 = 32'd72; 
32'd478: dataIn2 = 32'd69; 
32'd479: dataIn2 = 32'd4; 
32'd480: dataIn2 = 32'd78; 
32'd481: dataIn2 = 32'd3; 
32'd482: dataIn2 = 32'd68; 
32'd483: dataIn2 = 32'd9; 
32'd484: dataIn2 = 32'd17; 
32'd485: dataIn2 = 32'd7; 
32'd486: dataIn2 = 32'd49; 
32'd487: dataIn2 = 32'd71; 
32'd488: dataIn2 = 32'd52; 
32'd489: dataIn2 = 32'd42; 
32'd490: dataIn2 = 32'd36; 
32'd491: dataIn2 = 32'd8; 
32'd492: dataIn2 = 32'd6; 
32'd493: dataIn2 = 32'd60; 
32'd494: dataIn2 = 32'd3; 
32'd495: dataIn2 = 32'd96; 
32'd496: dataIn2 = 32'd65; 
32'd497: dataIn2 = 32'd51; 
32'd498: dataIn2 = 32'd78; 
32'd499: dataIn2 = 32'd19; 
32'd500: dataIn2 = 32'd0; 
32'd501: dataIn2 = 32'd66; 
32'd502: dataIn2 = 32'd54; 
32'd503: dataIn2 = 32'd81; 
32'd504: dataIn2 = 32'd51; 
32'd505: dataIn2 = 32'd19; 
32'd506: dataIn2 = 32'd66; 
32'd507: dataIn2 = 32'd63; 
32'd508: dataIn2 = 32'd25; 
32'd509: dataIn2 = 32'd11; 
32'd510: dataIn2 = 32'd35; 
32'd511: dataIn2 = 32'd29; 
32'd512: dataIn2 = 32'd41; 
32'd513: dataIn2 = 32'd55; 
32'd514: dataIn2 = 32'd63; 
32'd515: dataIn2 = 32'd15; 
32'd516: dataIn2 = 32'd74; 
32'd517: dataIn2 = 32'd30; 
32'd518: dataIn2 = 32'd75; 
32'd519: dataIn2 = 32'd40; 
32'd520: dataIn2 = 32'd6; 
32'd521: dataIn2 = 32'd17; 
32'd522: dataIn2 = 32'd87; 
32'd523: dataIn2 = 32'd18; 
32'd524: dataIn2 = 32'd10; 
32'd525: dataIn2 = 32'd37; 
32'd526: dataIn2 = 32'd81; 
32'd527: dataIn2 = 32'd60; 
32'd528: dataIn2 = 32'd25; 
32'd529: dataIn2 = 32'd6; 
32'd530: dataIn2 = 32'd27; 
32'd531: dataIn2 = 32'd82; 
32'd532: dataIn2 = 32'd98; 
32'd533: dataIn2 = 32'd2; 
32'd534: dataIn2 = 32'd96; 
32'd535: dataIn2 = 32'd59; 
32'd536: dataIn2 = 32'd78; 
32'd537: dataIn2 = 32'd20; 
32'd538: dataIn2 = 32'd18; 
32'd539: dataIn2 = 32'd99; 
32'd540: dataIn2 = 32'd30; 
32'd541: dataIn2 = 32'd56; 
32'd542: dataIn2 = 32'd0; 
32'd543: dataIn2 = 32'd25; 
32'd544: dataIn2 = 32'd29; 
32'd545: dataIn2 = 32'd54; 
32'd546: dataIn2 = 32'd34; 
32'd547: dataIn2 = 32'd48; 
32'd548: dataIn2 = 32'd34; 
32'd549: dataIn2 = 32'd44; 
32'd550: dataIn2 = 32'd82; 
32'd551: dataIn2 = 32'd89; 
32'd552: dataIn2 = 32'd89; 
32'd553: dataIn2 = 32'd87; 
32'd554: dataIn2 = 32'd26; 
32'd555: dataIn2 = 32'd18; 
32'd556: dataIn2 = 32'd53; 
32'd557: dataIn2 = 32'd23; 
32'd558: dataIn2 = 32'd10; 
32'd559: dataIn2 = 32'd8; 
32'd560: dataIn2 = 32'd30; 
32'd561: dataIn2 = 32'd2; 
32'd562: dataIn2 = 32'd71; 
32'd563: dataIn2 = 32'd11; 
32'd564: dataIn2 = 32'd14; 
32'd565: dataIn2 = 32'd80; 
32'd566: dataIn2 = 32'd94; 
32'd567: dataIn2 = 32'd20; 
32'd568: dataIn2 = 32'd94; 
32'd569: dataIn2 = 32'd13; 
32'd570: dataIn2 = 32'd7; 
32'd571: dataIn2 = 32'd98; 
32'd572: dataIn2 = 32'd61; 
32'd573: dataIn2 = 32'd82; 
32'd574: dataIn2 = 32'd71; 
32'd575: dataIn2 = 32'd24; 
32'd576: dataIn2 = 32'd36; 
32'd577: dataIn2 = 32'd36; 
32'd578: dataIn2 = 32'd96; 
32'd579: dataIn2 = 32'd100; 
32'd580: dataIn2 = 32'd43; 
32'd581: dataIn2 = 32'd14; 
32'd582: dataIn2 = 32'd75; 
32'd583: dataIn2 = 32'd77; 
32'd584: dataIn2 = 32'd90; 
32'd585: dataIn2 = 32'd3; 
32'd586: dataIn2 = 32'd7; 
32'd587: dataIn2 = 32'd93; 
32'd588: dataIn2 = 32'd81; 
32'd589: dataIn2 = 32'd30; 
32'd590: dataIn2 = 32'd10; 
32'd591: dataIn2 = 32'd50; 
32'd592: dataIn2 = 32'd89; 
32'd593: dataIn2 = 32'd91; 
32'd594: dataIn2 = 32'd84; 
32'd595: dataIn2 = 32'd29; 
32'd596: dataIn2 = 32'd7; 
32'd597: dataIn2 = 32'd19; 
32'd598: dataIn2 = 32'd78; 
32'd599: dataIn2 = 32'd17; 
32'd600: dataIn2 = 32'd0; 
32'd601: dataIn2 = 32'd86; 
32'd602: dataIn2 = 32'd39; 
32'd603: dataIn2 = 32'd60; 
32'd604: dataIn2 = 32'd15; 
32'd605: dataIn2 = 32'd17; 
32'd606: dataIn2 = 32'd54; 
32'd607: dataIn2 = 32'd69; 
32'd608: dataIn2 = 32'd40; 
32'd609: dataIn2 = 32'd33; 
32'd610: dataIn2 = 32'd69; 
32'd611: dataIn2 = 32'd57; 
32'd612: dataIn2 = 32'd15; 
32'd613: dataIn2 = 32'd27; 
32'd614: dataIn2 = 32'd15; 
32'd615: dataIn2 = 32'd72; 
32'd616: dataIn2 = 32'd69; 
32'd617: dataIn2 = 32'd55; 
32'd618: dataIn2 = 32'd26; 
32'd619: dataIn2 = 32'd54; 
32'd620: dataIn2 = 32'd22; 
32'd621: dataIn2 = 32'd11; 
32'd622: dataIn2 = 32'd38; 
32'd623: dataIn2 = 32'd24; 
32'd624: dataIn2 = 32'd52; 
32'd625: dataIn2 = 32'd9; 
32'd626: dataIn2 = 32'd56; 
32'd627: dataIn2 = 32'd38; 
32'd628: dataIn2 = 32'd66; 
32'd629: dataIn2 = 32'd73; 
32'd630: dataIn2 = 32'd97; 
32'd631: dataIn2 = 32'd66; 
32'd632: dataIn2 = 32'd1; 
32'd633: dataIn2 = 32'd88; 
32'd634: dataIn2 = 32'd50; 
32'd635: dataIn2 = 32'd24; 
32'd636: dataIn2 = 32'd39; 
32'd637: dataIn2 = 32'd93; 
32'd638: dataIn2 = 32'd77; 
32'd639: dataIn2 = 32'd38; 
32'd640: dataIn2 = 32'd98; 
32'd641: dataIn2 = 32'd81; 
32'd642: dataIn2 = 32'd50; 
32'd643: dataIn2 = 32'd71; 
32'd644: dataIn2 = 32'd23; 
32'd645: dataIn2 = 32'd91; 
32'd646: dataIn2 = 32'd38; 
32'd647: dataIn2 = 32'd8; 
32'd648: dataIn2 = 32'd87; 
32'd649: dataIn2 = 32'd42; 
32'd650: dataIn2 = 32'd100; 
32'd651: dataIn2 = 32'd59; 
32'd652: dataIn2 = 32'd19; 
32'd653: dataIn2 = 32'd77; 
32'd654: dataIn2 = 32'd71; 
32'd655: dataIn2 = 32'd84; 
32'd656: dataIn2 = 32'd79; 
32'd657: dataIn2 = 32'd47; 
32'd658: dataIn2 = 32'd17; 
32'd659: dataIn2 = 32'd53; 
32'd660: dataIn2 = 32'd22; 
32'd661: dataIn2 = 32'd4; 
32'd662: dataIn2 = 32'd84; 
32'd663: dataIn2 = 32'd11; 
32'd664: dataIn2 = 32'd5; 
32'd665: dataIn2 = 32'd75; 
32'd666: dataIn2 = 32'd71; 
32'd667: dataIn2 = 32'd1; 
32'd668: dataIn2 = 32'd99; 
32'd669: dataIn2 = 32'd23; 
32'd670: dataIn2 = 32'd18; 
32'd671: dataIn2 = 32'd73; 
32'd672: dataIn2 = 32'd42; 
32'd673: dataIn2 = 32'd87; 
32'd674: dataIn2 = 32'd22; 
32'd675: dataIn2 = 32'd84; 
32'd676: dataIn2 = 32'd56; 
32'd677: dataIn2 = 32'd61; 
32'd678: dataIn2 = 32'd96; 
32'd679: dataIn2 = 32'd87; 
32'd680: dataIn2 = 32'd98; 
32'd681: dataIn2 = 32'd13; 
32'd682: dataIn2 = 32'd11; 
32'd683: dataIn2 = 32'd11; 
32'd684: dataIn2 = 32'd41; 
32'd685: dataIn2 = 32'd48; 
32'd686: dataIn2 = 32'd85; 
32'd687: dataIn2 = 32'd28; 
32'd688: dataIn2 = 32'd68; 
32'd689: dataIn2 = 32'd49; 
32'd690: dataIn2 = 32'd65; 
32'd691: dataIn2 = 32'd5; 
32'd692: dataIn2 = 32'd31; 
32'd693: dataIn2 = 32'd7; 
32'd694: dataIn2 = 32'd15; 
32'd695: dataIn2 = 32'd59; 
32'd696: dataIn2 = 32'd11; 
32'd697: dataIn2 = 32'd58; 
32'd698: dataIn2 = 32'd60; 
32'd699: dataIn2 = 32'd62; 
32'd700: dataIn2 = 32'd63; 
32'd701: dataIn2 = 32'd36; 
32'd702: dataIn2 = 32'd72; 
32'd703: dataIn2 = 32'd42; 
32'd704: dataIn2 = 32'd64; 
32'd705: dataIn2 = 32'd43; 
32'd706: dataIn2 = 32'd22; 
32'd707: dataIn2 = 32'd66; 
32'd708: dataIn2 = 32'd71; 
32'd709: dataIn2 = 32'd37; 
32'd710: dataIn2 = 32'd93; 
32'd711: dataIn2 = 32'd79; 
32'd712: dataIn2 = 32'd16; 
32'd713: dataIn2 = 32'd29; 
32'd714: dataIn2 = 32'd75; 
32'd715: dataIn2 = 32'd1; 
32'd716: dataIn2 = 32'd64; 
32'd717: dataIn2 = 32'd73; 
32'd718: dataIn2 = 32'd86; 
32'd719: dataIn2 = 32'd57; 
32'd720: dataIn2 = 32'd64; 
32'd721: dataIn2 = 32'd33; 
32'd722: dataIn2 = 32'd4; 
32'd723: dataIn2 = 32'd74; 
32'd724: dataIn2 = 32'd2; 
32'd725: dataIn2 = 32'd27; 
32'd726: dataIn2 = 32'd89; 
32'd727: dataIn2 = 32'd67; 
32'd728: dataIn2 = 32'd69; 
32'd729: dataIn2 = 32'd62; 
32'd730: dataIn2 = 32'd11; 
32'd731: dataIn2 = 32'd10; 
32'd732: dataIn2 = 32'd85; 
32'd733: dataIn2 = 32'd30; 
32'd734: dataIn2 = 32'd25; 
32'd735: dataIn2 = 32'd55; 
32'd736: dataIn2 = 32'd94; 
32'd737: dataIn2 = 32'd80; 
32'd738: dataIn2 = 32'd24; 
32'd739: dataIn2 = 32'd80; 
32'd740: dataIn2 = 32'd15; 
32'd741: dataIn2 = 32'd77; 
32'd742: dataIn2 = 32'd1; 
32'd743: dataIn2 = 32'd20; 
32'd744: dataIn2 = 32'd37; 
32'd745: dataIn2 = 32'd18; 
32'd746: dataIn2 = 32'd62; 
32'd747: dataIn2 = 32'd82; 
32'd748: dataIn2 = 32'd57; 
32'd749: dataIn2 = 32'd89; 
32'd750: dataIn2 = 32'd36; 
32'd751: dataIn2 = 32'd80; 
32'd752: dataIn2 = 32'd67; 
32'd753: dataIn2 = 32'd5; 
32'd754: dataIn2 = 32'd85; 
32'd755: dataIn2 = 32'd2; 
32'd756: dataIn2 = 32'd74; 
32'd757: dataIn2 = 32'd24; 
32'd758: dataIn2 = 32'd74; 
32'd759: dataIn2 = 32'd78; 
32'd760: dataIn2 = 32'd22; 
32'd761: dataIn2 = 32'd54; 
32'd762: dataIn2 = 32'd93; 
32'd763: dataIn2 = 32'd43; 
32'd764: dataIn2 = 32'd93; 
32'd765: dataIn2 = 32'd2; 
32'd766: dataIn2 = 32'd47; 
32'd767: dataIn2 = 32'd13; 
32'd768: dataIn2 = 32'd84; 
32'd769: dataIn2 = 32'd59; 
32'd770: dataIn2 = 32'd90; 
32'd771: dataIn2 = 32'd78; 
32'd772: dataIn2 = 32'd85; 
32'd773: dataIn2 = 32'd39; 
32'd774: dataIn2 = 32'd71; 
32'd775: dataIn2 = 32'd74; 
32'd776: dataIn2 = 32'd99; 
32'd777: dataIn2 = 32'd28; 
32'd778: dataIn2 = 32'd69; 
32'd779: dataIn2 = 32'd33; 
32'd780: dataIn2 = 32'd84; 
32'd781: dataIn2 = 32'd36; 
32'd782: dataIn2 = 32'd52; 
32'd783: dataIn2 = 32'd74; 
32'd784: dataIn2 = 32'd18; 
32'd785: dataIn2 = 32'd10; 
32'd786: dataIn2 = 32'd60; 
32'd787: dataIn2 = 32'd68; 
32'd788: dataIn2 = 32'd22; 
32'd789: dataIn2 = 32'd67; 
32'd790: dataIn2 = 32'd1; 
32'd791: dataIn2 = 32'd91; 
32'd792: dataIn2 = 32'd29; 
32'd793: dataIn2 = 32'd8; 
32'd794: dataIn2 = 32'd37; 
32'd795: dataIn2 = 32'd76; 
32'd796: dataIn2 = 32'd7; 
32'd797: dataIn2 = 32'd27; 
32'd798: dataIn2 = 32'd54; 
32'd799: dataIn2 = 32'd67; 
32'd800: dataIn2 = 32'd61; 
32'd801: dataIn2 = 32'd91; 
32'd802: dataIn2 = 32'd37; 
32'd803: dataIn2 = 32'd47; 
32'd804: dataIn2 = 32'd8; 
32'd805: dataIn2 = 32'd45; 
32'd806: dataIn2 = 32'd39; 
32'd807: dataIn2 = 32'd3; 
32'd808: dataIn2 = 32'd50; 
32'd809: dataIn2 = 32'd18; 
32'd810: dataIn2 = 32'd100; 
32'd811: dataIn2 = 32'd64; 
32'd812: dataIn2 = 32'd27; 
32'd813: dataIn2 = 32'd43; 
32'd814: dataIn2 = 32'd50; 
32'd815: dataIn2 = 32'd7; 
32'd816: dataIn2 = 32'd68; 
32'd817: dataIn2 = 32'd72; 
32'd818: dataIn2 = 32'd47; 
32'd819: dataIn2 = 32'd30; 
32'd820: dataIn2 = 32'd19; 
32'd821: dataIn2 = 32'd76; 
32'd822: dataIn2 = 32'd4; 
32'd823: dataIn2 = 32'd12; 
32'd824: dataIn2 = 32'd38; 
32'd825: dataIn2 = 32'd15; 
32'd826: dataIn2 = 32'd2; 
32'd827: dataIn2 = 32'd71; 
32'd828: dataIn2 = 32'd12; 
32'd829: dataIn2 = 32'd26; 
32'd830: dataIn2 = 32'd73; 
32'd831: dataIn2 = 32'd41; 
32'd832: dataIn2 = 32'd51; 
32'd833: dataIn2 = 32'd7; 
32'd834: dataIn2 = 32'd97; 
32'd835: dataIn2 = 32'd80; 
32'd836: dataIn2 = 32'd71; 
32'd837: dataIn2 = 32'd89; 
32'd838: dataIn2 = 32'd88; 
32'd839: dataIn2 = 32'd53; 
32'd840: dataIn2 = 32'd94; 
32'd841: dataIn2 = 32'd61; 
32'd842: dataIn2 = 32'd31; 
32'd843: dataIn2 = 32'd87; 
32'd844: dataIn2 = 32'd59; 
32'd845: dataIn2 = 32'd83; 
32'd846: dataIn2 = 32'd10; 
32'd847: dataIn2 = 32'd31; 
32'd848: dataIn2 = 32'd87; 
32'd849: dataIn2 = 32'd30; 
32'd850: dataIn2 = 32'd85; 
32'd851: dataIn2 = 32'd70; 
32'd852: dataIn2 = 32'd75; 
32'd853: dataIn2 = 32'd7; 
32'd854: dataIn2 = 32'd85; 
32'd855: dataIn2 = 32'd84; 
32'd856: dataIn2 = 32'd56; 
32'd857: dataIn2 = 32'd45; 
32'd858: dataIn2 = 32'd3; 
32'd859: dataIn2 = 32'd78; 
32'd860: dataIn2 = 32'd28; 
32'd861: dataIn2 = 32'd74; 
32'd862: dataIn2 = 32'd75; 
32'd863: dataIn2 = 32'd29; 
32'd864: dataIn2 = 32'd94; 
32'd865: dataIn2 = 32'd12; 
32'd866: dataIn2 = 32'd58; 
32'd867: dataIn2 = 32'd44; 
32'd868: dataIn2 = 32'd70; 
32'd869: dataIn2 = 32'd39; 
32'd870: dataIn2 = 32'd73; 
32'd871: dataIn2 = 32'd8; 
32'd872: dataIn2 = 32'd24; 
32'd873: dataIn2 = 32'd76; 
32'd874: dataIn2 = 32'd60; 
32'd875: dataIn2 = 32'd95; 
32'd876: dataIn2 = 32'd18; 
32'd877: dataIn2 = 32'd91; 
32'd878: dataIn2 = 32'd36; 
32'd879: dataIn2 = 32'd1; 
32'd880: dataIn2 = 32'd37; 
32'd881: dataIn2 = 32'd97; 
32'd882: dataIn2 = 32'd45; 
32'd883: dataIn2 = 32'd80; 
32'd884: dataIn2 = 32'd59; 
32'd885: dataIn2 = 32'd3; 
32'd886: dataIn2 = 32'd92; 
32'd887: dataIn2 = 32'd40; 
32'd888: dataIn2 = 32'd17; 
32'd889: dataIn2 = 32'd36; 
32'd890: dataIn2 = 32'd44; 
32'd891: dataIn2 = 32'd28; 
32'd892: dataIn2 = 32'd17; 
32'd893: dataIn2 = 32'd51; 
32'd894: dataIn2 = 32'd8; 
32'd895: dataIn2 = 32'd92; 
32'd896: dataIn2 = 32'd48; 
32'd897: dataIn2 = 32'd55; 
32'd898: dataIn2 = 32'd13; 
32'd899: dataIn2 = 32'd84; 
32'd900: dataIn2 = 32'd27; 
32'd901: dataIn2 = 32'd28; 
32'd902: dataIn2 = 32'd89; 
32'd903: dataIn2 = 32'd18; 
32'd904: dataIn2 = 32'd8; 
32'd905: dataIn2 = 32'd61; 
32'd906: dataIn2 = 32'd51; 
32'd907: dataIn2 = 32'd41; 
32'd908: dataIn2 = 32'd36; 
32'd909: dataIn2 = 32'd47; 
32'd910: dataIn2 = 32'd26; 
32'd911: dataIn2 = 32'd51; 
32'd912: dataIn2 = 32'd84; 
32'd913: dataIn2 = 32'd24; 
32'd914: dataIn2 = 32'd29; 
32'd915: dataIn2 = 32'd33; 
32'd916: dataIn2 = 32'd8; 
32'd917: dataIn2 = 32'd23; 
32'd918: dataIn2 = 32'd98; 
32'd919: dataIn2 = 32'd3; 
32'd920: dataIn2 = 32'd68; 
32'd921: dataIn2 = 32'd93; 
32'd922: dataIn2 = 32'd76; 
32'd923: dataIn2 = 32'd61; 
32'd924: dataIn2 = 32'd27; 
32'd925: dataIn2 = 32'd6; 
32'd926: dataIn2 = 32'd77; 
32'd927: dataIn2 = 32'd74; 
32'd928: dataIn2 = 32'd18; 
32'd929: dataIn2 = 32'd83; 
32'd930: dataIn2 = 32'd85; 
32'd931: dataIn2 = 32'd22; 
32'd932: dataIn2 = 32'd38; 
32'd933: dataIn2 = 32'd47; 
32'd934: dataIn2 = 32'd92; 
32'd935: dataIn2 = 32'd28; 
32'd936: dataIn2 = 32'd78; 
32'd937: dataIn2 = 32'd2; 
32'd938: dataIn2 = 32'd98; 
32'd939: dataIn2 = 32'd72; 
32'd940: dataIn2 = 32'd36; 
32'd941: dataIn2 = 32'd74; 
32'd942: dataIn2 = 32'd4; 
32'd943: dataIn2 = 32'd25; 
32'd944: dataIn2 = 32'd42; 
32'd945: dataIn2 = 32'd60; 
32'd946: dataIn2 = 32'd70; 
32'd947: dataIn2 = 32'd44; 
32'd948: dataIn2 = 32'd66; 
32'd949: dataIn2 = 32'd52; 
32'd950: dataIn2 = 32'd89; 
32'd951: dataIn2 = 32'd57; 
32'd952: dataIn2 = 32'd68; 
32'd953: dataIn2 = 32'd21; 
32'd954: dataIn2 = 32'd67; 
32'd955: dataIn2 = 32'd31; 
32'd956: dataIn2 = 32'd60; 
32'd957: dataIn2 = 32'd12; 
32'd958: dataIn2 = 32'd3; 
32'd959: dataIn2 = 32'd25; 
32'd960: dataIn2 = 32'd15; 
32'd961: dataIn2 = 32'd27; 
32'd962: dataIn2 = 32'd51; 
32'd963: dataIn2 = 32'd26; 
32'd964: dataIn2 = 32'd41; 
32'd965: dataIn2 = 32'd9; 
32'd966: dataIn2 = 32'd48; 
32'd967: dataIn2 = 32'd51; 
32'd968: dataIn2 = 32'd66; 
32'd969: dataIn2 = 32'd10; 
32'd970: dataIn2 = 32'd17; 
32'd971: dataIn2 = 32'd81; 
32'd972: dataIn2 = 32'd4; 
32'd973: dataIn2 = 32'd81; 
32'd974: dataIn2 = 32'd5; 
32'd975: dataIn2 = 32'd17; 
32'd976: dataIn2 = 32'd93; 
32'd977: dataIn2 = 32'd21; 
32'd978: dataIn2 = 32'd22; 
32'd979: dataIn2 = 32'd64; 
32'd980: dataIn2 = 32'd72; 
32'd981: dataIn2 = 32'd83; 
32'd982: dataIn2 = 32'd14; 
32'd983: dataIn2 = 32'd26; 
32'd984: dataIn2 = 32'd45; 
32'd985: dataIn2 = 32'd33; 
32'd986: dataIn2 = 32'd64; 
32'd987: dataIn2 = 32'd14; 
32'd988: dataIn2 = 32'd85; 
32'd989: dataIn2 = 32'd4; 
32'd990: dataIn2 = 32'd48; 
32'd991: dataIn2 = 32'd17; 
32'd992: dataIn2 = 32'd92; 
32'd993: dataIn2 = 32'd19; 
32'd994: dataIn2 = 32'd22; 
32'd995: dataIn2 = 32'd98; 
32'd996: dataIn2 = 32'd79; 
32'd997: dataIn2 = 32'd65; 
32'd998: dataIn2 = 32'd87; 
32'd999: dataIn2 = 32'd26; 
32'd1000: dataIn2 = 32'd24; 
32'd1001: dataIn2 = 32'd98; 
32'd1002: dataIn2 = 32'd90; 
32'd1003: dataIn2 = 32'd75; 
32'd1004: dataIn2 = 32'd54; 
32'd1005: dataIn2 = 32'd84; 
32'd1006: dataIn2 = 32'd72; 
32'd1007: dataIn2 = 32'd51; 
32'd1008: dataIn2 = 32'd59; 
32'd1009: dataIn2 = 32'd34; 
32'd1010: dataIn2 = 32'd49; 
32'd1011: dataIn2 = 32'd36; 
32'd1012: dataIn2 = 32'd27; 
32'd1013: dataIn2 = 32'd18; 
32'd1014: dataIn2 = 32'd18; 
32'd1015: dataIn2 = 32'd11; 
32'd1016: dataIn2 = 32'd37; 
32'd1017: dataIn2 = 32'd68; 
32'd1018: dataIn2 = 32'd68; 
32'd1019: dataIn2 = 32'd8; 
32'd1020: dataIn2 = 32'd25; 
32'd1021: dataIn2 = 32'd0; 
32'd1022: dataIn2 = 32'd64; 
32'd1023: dataIn2 = 32'd32; 
32'd1024: dataIn2 = 32'd19; 
32'd1025: dataIn2 = 32'd77; 
32'd1026: dataIn2 = 32'd96; 
32'd1027: dataIn2 = 32'd64; 
32'd1028: dataIn2 = 32'd0; 
32'd1029: dataIn2 = 32'd58; 
32'd1030: dataIn2 = 32'd74; 
32'd1031: dataIn2 = 32'd84; 
32'd1032: dataIn2 = 32'd63; 
32'd1033: dataIn2 = 32'd33; 
32'd1034: dataIn2 = 32'd14; 
32'd1035: dataIn2 = 32'd20; 
32'd1036: dataIn2 = 32'd44; 
32'd1037: dataIn2 = 32'd94; 
32'd1038: dataIn2 = 32'd78; 
32'd1039: dataIn2 = 32'd22; 
32'd1040: dataIn2 = 32'd99; 
32'd1041: dataIn2 = 32'd37; 
32'd1042: dataIn2 = 32'd37; 
32'd1043: dataIn2 = 32'd10; 
32'd1044: dataIn2 = 32'd77; 
32'd1045: dataIn2 = 32'd42; 
32'd1046: dataIn2 = 32'd83; 
32'd1047: dataIn2 = 32'd56; 
32'd1048: dataIn2 = 32'd62; 
32'd1049: dataIn2 = 32'd61; 
32'd1050: dataIn2 = 32'd1; 
32'd1051: dataIn2 = 32'd31; 
32'd1052: dataIn2 = 32'd74; 
32'd1053: dataIn2 = 32'd10; 
32'd1054: dataIn2 = 32'd23; 
32'd1055: dataIn2 = 32'd96; 
32'd1056: dataIn2 = 32'd90; 
32'd1057: dataIn2 = 32'd21; 
32'd1058: dataIn2 = 32'd57; 
32'd1059: dataIn2 = 32'd12; 
32'd1060: dataIn2 = 32'd31; 
32'd1061: dataIn2 = 32'd93; 
32'd1062: dataIn2 = 32'd60; 
32'd1063: dataIn2 = 32'd2; 
32'd1064: dataIn2 = 32'd53; 
32'd1065: dataIn2 = 32'd20; 
32'd1066: dataIn2 = 32'd43; 
32'd1067: dataIn2 = 32'd72; 
32'd1068: dataIn2 = 32'd68; 
32'd1069: dataIn2 = 32'd82; 
32'd1070: dataIn2 = 32'd62; 
32'd1071: dataIn2 = 32'd72; 
32'd1072: dataIn2 = 32'd71; 
32'd1073: dataIn2 = 32'd27; 
32'd1074: dataIn2 = 32'd60; 
32'd1075: dataIn2 = 32'd60; 
32'd1076: dataIn2 = 32'd49; 
32'd1077: dataIn2 = 32'd79; 
32'd1078: dataIn2 = 32'd10; 
32'd1079: dataIn2 = 32'd62; 
32'd1080: dataIn2 = 32'd21; 
32'd1081: dataIn2 = 32'd21; 
32'd1082: dataIn2 = 32'd58; 
32'd1083: dataIn2 = 32'd19; 
32'd1084: dataIn2 = 32'd43; 
32'd1085: dataIn2 = 32'd41; 
32'd1086: dataIn2 = 32'd36; 
32'd1087: dataIn2 = 32'd78; 
32'd1088: dataIn2 = 32'd33; 
32'd1089: dataIn2 = 32'd40; 
32'd1090: dataIn2 = 32'd43; 
32'd1091: dataIn2 = 32'd11; 
32'd1092: dataIn2 = 32'd32; 
32'd1093: dataIn2 = 32'd0; 
32'd1094: dataIn2 = 32'd11; 
32'd1095: dataIn2 = 32'd1; 
32'd1096: dataIn2 = 32'd60; 
32'd1097: dataIn2 = 32'd69; 
32'd1098: dataIn2 = 32'd82; 
32'd1099: dataIn2 = 32'd69; 
32'd1100: dataIn2 = 32'd100; 
32'd1101: dataIn2 = 32'd87; 
32'd1102: dataIn2 = 32'd20; 
32'd1103: dataIn2 = 32'd74; 
32'd1104: dataIn2 = 32'd4; 
32'd1105: dataIn2 = 32'd35; 
32'd1106: dataIn2 = 32'd32; 
32'd1107: dataIn2 = 32'd40; 
32'd1108: dataIn2 = 32'd19; 
32'd1109: dataIn2 = 32'd9; 
32'd1110: dataIn2 = 32'd3; 
32'd1111: dataIn2 = 32'd16; 
32'd1112: dataIn2 = 32'd85; 
32'd1113: dataIn2 = 32'd59; 
32'd1114: dataIn2 = 32'd70; 
32'd1115: dataIn2 = 32'd50; 
32'd1116: dataIn2 = 32'd80; 
32'd1117: dataIn2 = 32'd46; 
32'd1118: dataIn2 = 32'd24; 
32'd1119: dataIn2 = 32'd2; 
32'd1120: dataIn2 = 32'd65; 
32'd1121: dataIn2 = 32'd14; 
32'd1122: dataIn2 = 32'd31; 
32'd1123: dataIn2 = 32'd15; 
32'd1124: dataIn2 = 32'd5; 
32'd1125: dataIn2 = 32'd27; 
32'd1126: dataIn2 = 32'd68; 
32'd1127: dataIn2 = 32'd66; 
32'd1128: dataIn2 = 32'd88; 
32'd1129: dataIn2 = 32'd58; 
32'd1130: dataIn2 = 32'd67; 
32'd1131: dataIn2 = 32'd84; 
32'd1132: dataIn2 = 32'd19; 
32'd1133: dataIn2 = 32'd52; 
32'd1134: dataIn2 = 32'd84; 
32'd1135: dataIn2 = 32'd14; 
32'd1136: dataIn2 = 32'd9; 
32'd1137: dataIn2 = 32'd54; 
32'd1138: dataIn2 = 32'd97; 
32'd1139: dataIn2 = 32'd32; 
32'd1140: dataIn2 = 32'd49; 
32'd1141: dataIn2 = 32'd70; 
32'd1142: dataIn2 = 32'd79; 
32'd1143: dataIn2 = 32'd27; 
32'd1144: dataIn2 = 32'd9; 
32'd1145: dataIn2 = 32'd77; 
32'd1146: dataIn2 = 32'd62; 
32'd1147: dataIn2 = 32'd69; 
32'd1148: dataIn2 = 32'd44; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_64_80.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
