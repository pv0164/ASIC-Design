//32x32 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 512 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
  wire [31:0]addr1,addr2; 
  wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base,row_base,matrix_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,v_values_base,wdata_col_base,matrix_base,addr1,addr2,dataIn1,dataIn2,Rst,row_base,RD,csize);  //frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  v_values_base = 32'd2; 
  matrix_base = 32'd170 ; 
  wdata_col_base = 32'd6820 ; 
  row_base = 32'd73320 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #10420; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd73320: dataIn1 = 32'd0
; 
32'd73321: dataIn1 = 32'd17
; 
32'd73322: dataIn1 = 32'd33
; 
32'd73323: dataIn1 = 32'd47
; 
32'd73324: dataIn1 = 32'd65
; 
32'd73325: dataIn1 = 32'd79
; 
32'd73326: dataIn1 = 32'd95
; 
32'd73327: dataIn1 = 32'd112
; 
32'd73328: dataIn1 = 32'd130
; 
32'd73329: dataIn1 = 32'd146
; 
32'd73330: dataIn1 = 32'd159
; 
32'd73331: dataIn1 = 32'd178
; 
32'd73332: dataIn1 = 32'd191
; 
32'd73333: dataIn1 = 32'd208
; 
32'd73334: dataIn1 = 32'd223
; 
32'd73335: dataIn1 = 32'd237
; 
32'd73336: dataIn1 = 32'd252
; 
32'd73337: dataIn1 = 32'd274
; 
32'd73338: dataIn1 = 32'd296
; 
32'd73339: dataIn1 = 32'd307
; 
32'd73340: dataIn1 = 32'd320
; 
32'd73341: dataIn1 = 32'd333
; 
32'd73342: dataIn1 = 32'd345
; 
32'd73343: dataIn1 = 32'd360
; 
32'd73344: dataIn1 = 32'd372
; 
32'd73345: dataIn1 = 32'd386
; 
32'd73346: dataIn1 = 32'd405
; 
32'd73347: dataIn1 = 32'd419
; 
32'd73348: dataIn1 = 32'd437
; 
32'd73349: dataIn1 = 32'd452
; 
32'd73350: dataIn1 = 32'd473
; 
32'd73351: dataIn1 = 32'd483
; 
32'd73352: dataIn1 = 32'd499
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
32'd6820: dataIn1 = 32'd0
; 
32'd6821: dataIn1 = 32'd17
; 
32'd6822: dataIn1 = 32'd33
; 
32'd6823: dataIn1 = 32'd47
; 
32'd6824: dataIn1 = 32'd65
; 
32'd6825: dataIn1 = 32'd79
; 
32'd6826: dataIn1 = 32'd95
; 
32'd6827: dataIn1 = 32'd112
; 
32'd6828: dataIn1 = 32'd130
; 
32'd6829: dataIn1 = 32'd146
; 
32'd6830: dataIn1 = 32'd159
; 
32'd6831: dataIn1 = 32'd178
; 
32'd6832: dataIn1 = 32'd191
; 
32'd6833: dataIn1 = 32'd208
; 
32'd6834: dataIn1 = 32'd223
; 
32'd6835: dataIn1 = 32'd237
; 
32'd6836: dataIn1 = 32'd252
; 
32'd6837: dataIn1 = 32'd274
; 
32'd6838: dataIn1 = 32'd296
; 
32'd6839: dataIn1 = 32'd307
; 
32'd6840: dataIn1 = 32'd320
; 
32'd6841: dataIn1 = 32'd333
; 
32'd6842: dataIn1 = 32'd345
; 
32'd6843: dataIn1 = 32'd360
; 
32'd6844: dataIn1 = 32'd372
; 
32'd6845: dataIn1 = 32'd386
; 
32'd6846: dataIn1 = 32'd405
; 
32'd6847: dataIn1 = 32'd419
; 
32'd6848: dataIn1 = 32'd437
; 
32'd6849: dataIn1 = 32'd452
; 
32'd6850: dataIn1 = 32'd473
; 
32'd6851: dataIn1 = 32'd483
; 
32'd6852: dataIn1 = 32'd499
; 
32'd6853: dataIn1 = 32'd1
; 
32'd6854: dataIn1 = 32'd2
; 
32'd6855: dataIn1 = 32'd3
; 
32'd6856: dataIn1 = 32'd5
; 
32'd6857: dataIn1 = 32'd12
; 
32'd6858: dataIn1 = 32'd13
; 
32'd6859: dataIn1 = 32'd14
; 
32'd6860: dataIn1 = 32'd16
; 
32'd6861: dataIn1 = 32'd18
; 
32'd6862: dataIn1 = 32'd19
; 
32'd6863: dataIn1 = 32'd20
; 
32'd6864: dataIn1 = 32'd21
; 
32'd6865: dataIn1 = 32'd23
; 
32'd6866: dataIn1 = 32'd28
; 
32'd6867: dataIn1 = 32'd29
; 
32'd6868: dataIn1 = 32'd30
; 
32'd6869: dataIn1 = 32'd31
; 
32'd6870: dataIn1 = 32'd0
; 
32'd6871: dataIn1 = 32'd2
; 
32'd6872: dataIn1 = 32'd4
; 
32'd6873: dataIn1 = 32'd5
; 
32'd6874: dataIn1 = 32'd10
; 
32'd6875: dataIn1 = 32'd11
; 
32'd6876: dataIn1 = 32'd12
; 
32'd6877: dataIn1 = 32'd14
; 
32'd6878: dataIn1 = 32'd17
; 
32'd6879: dataIn1 = 32'd20
; 
32'd6880: dataIn1 = 32'd21
; 
32'd6881: dataIn1 = 32'd22
; 
32'd6882: dataIn1 = 32'd25
; 
32'd6883: dataIn1 = 32'd26
; 
32'd6884: dataIn1 = 32'd28
; 
32'd6885: dataIn1 = 32'd31
; 
32'd6886: dataIn1 = 32'd2
; 
32'd6887: dataIn1 = 32'd6
; 
32'd6888: dataIn1 = 32'd7
; 
32'd6889: dataIn1 = 32'd10
; 
32'd6890: dataIn1 = 32'd11
; 
32'd6891: dataIn1 = 32'd13
; 
32'd6892: dataIn1 = 32'd16
; 
32'd6893: dataIn1 = 32'd17
; 
32'd6894: dataIn1 = 32'd18
; 
32'd6895: dataIn1 = 32'd22
; 
32'd6896: dataIn1 = 32'd24
; 
32'd6897: dataIn1 = 32'd29
; 
32'd6898: dataIn1 = 32'd30
; 
32'd6899: dataIn1 = 32'd31
; 
32'd6900: dataIn1 = 32'd0
; 
32'd6901: dataIn1 = 32'd2
; 
32'd6902: dataIn1 = 32'd3
; 
32'd6903: dataIn1 = 32'd5
; 
32'd6904: dataIn1 = 32'd6
; 
32'd6905: dataIn1 = 32'd8
; 
32'd6906: dataIn1 = 32'd9
; 
32'd6907: dataIn1 = 32'd10
; 
32'd6908: dataIn1 = 32'd11
; 
32'd6909: dataIn1 = 32'd12
; 
32'd6910: dataIn1 = 32'd13
; 
32'd6911: dataIn1 = 32'd15
; 
32'd6912: dataIn1 = 32'd18
; 
32'd6913: dataIn1 = 32'd20
; 
32'd6914: dataIn1 = 32'd23
; 
32'd6915: dataIn1 = 32'd25
; 
32'd6916: dataIn1 = 32'd27
; 
32'd6917: dataIn1 = 32'd28
; 
32'd6918: dataIn1 = 32'd4
; 
32'd6919: dataIn1 = 32'd5
; 
32'd6920: dataIn1 = 32'd7
; 
32'd6921: dataIn1 = 32'd8
; 
32'd6922: dataIn1 = 32'd9
; 
32'd6923: dataIn1 = 32'd11
; 
32'd6924: dataIn1 = 32'd14
; 
32'd6925: dataIn1 = 32'd17
; 
32'd6926: dataIn1 = 32'd19
; 
32'd6927: dataIn1 = 32'd22
; 
32'd6928: dataIn1 = 32'd23
; 
32'd6929: dataIn1 = 32'd24
; 
32'd6930: dataIn1 = 32'd26
; 
32'd6931: dataIn1 = 32'd31
; 
32'd6932: dataIn1 = 32'd1
; 
32'd6933: dataIn1 = 32'd2
; 
32'd6934: dataIn1 = 32'd4
; 
32'd6935: dataIn1 = 32'd5
; 
32'd6936: dataIn1 = 32'd6
; 
32'd6937: dataIn1 = 32'd7
; 
32'd6938: dataIn1 = 32'd12
; 
32'd6939: dataIn1 = 32'd13
; 
32'd6940: dataIn1 = 32'd15
; 
32'd6941: dataIn1 = 32'd16
; 
32'd6942: dataIn1 = 32'd19
; 
32'd6943: dataIn1 = 32'd23
; 
32'd6944: dataIn1 = 32'd25
; 
32'd6945: dataIn1 = 32'd26
; 
32'd6946: dataIn1 = 32'd27
; 
32'd6947: dataIn1 = 32'd29
; 
32'd6948: dataIn1 = 32'd1
; 
32'd6949: dataIn1 = 32'd3
; 
32'd6950: dataIn1 = 32'd9
; 
32'd6951: dataIn1 = 32'd10
; 
32'd6952: dataIn1 = 32'd11
; 
32'd6953: dataIn1 = 32'd12
; 
32'd6954: dataIn1 = 32'd13
; 
32'd6955: dataIn1 = 32'd16
; 
32'd6956: dataIn1 = 32'd18
; 
32'd6957: dataIn1 = 32'd20
; 
32'd6958: dataIn1 = 32'd21
; 
32'd6959: dataIn1 = 32'd22
; 
32'd6960: dataIn1 = 32'd23
; 
32'd6961: dataIn1 = 32'd26
; 
32'd6962: dataIn1 = 32'd27
; 
32'd6963: dataIn1 = 32'd30
; 
32'd6964: dataIn1 = 32'd31
; 
32'd6965: dataIn1 = 32'd0
; 
32'd6966: dataIn1 = 32'd1
; 
32'd6967: dataIn1 = 32'd2
; 
32'd6968: dataIn1 = 32'd3
; 
32'd6969: dataIn1 = 32'd4
; 
32'd6970: dataIn1 = 32'd7
; 
32'd6971: dataIn1 = 32'd13
; 
32'd6972: dataIn1 = 32'd15
; 
32'd6973: dataIn1 = 32'd16
; 
32'd6974: dataIn1 = 32'd17
; 
32'd6975: dataIn1 = 32'd18
; 
32'd6976: dataIn1 = 32'd20
; 
32'd6977: dataIn1 = 32'd22
; 
32'd6978: dataIn1 = 32'd25
; 
32'd6979: dataIn1 = 32'd26
; 
32'd6980: dataIn1 = 32'd27
; 
32'd6981: dataIn1 = 32'd29
; 
32'd6982: dataIn1 = 32'd31
; 
32'd6983: dataIn1 = 32'd1
; 
32'd6984: dataIn1 = 32'd2
; 
32'd6985: dataIn1 = 32'd3
; 
32'd6986: dataIn1 = 32'd4
; 
32'd6987: dataIn1 = 32'd8
; 
32'd6988: dataIn1 = 32'd10
; 
32'd6989: dataIn1 = 32'd11
; 
32'd6990: dataIn1 = 32'd12
; 
32'd6991: dataIn1 = 32'd14
; 
32'd6992: dataIn1 = 32'd21
; 
32'd6993: dataIn1 = 32'd22
; 
32'd6994: dataIn1 = 32'd24
; 
32'd6995: dataIn1 = 32'd26
; 
32'd6996: dataIn1 = 32'd27
; 
32'd6997: dataIn1 = 32'd28
; 
32'd6998: dataIn1 = 32'd31
; 
32'd6999: dataIn1 = 32'd0
; 
32'd7000: dataIn1 = 32'd6
; 
32'd7001: dataIn1 = 32'd7
; 
32'd7002: dataIn1 = 32'd8
; 
32'd7003: dataIn1 = 32'd9
; 
32'd7004: dataIn1 = 32'd10
; 
32'd7005: dataIn1 = 32'd14
; 
32'd7006: dataIn1 = 32'd18
; 
32'd7007: dataIn1 = 32'd20
; 
32'd7008: dataIn1 = 32'd21
; 
32'd7009: dataIn1 = 32'd23
; 
32'd7010: dataIn1 = 32'd27
; 
32'd7011: dataIn1 = 32'd31
; 
32'd7012: dataIn1 = 32'd0
; 
32'd7013: dataIn1 = 32'd3
; 
32'd7014: dataIn1 = 32'd4
; 
32'd7015: dataIn1 = 32'd5
; 
32'd7016: dataIn1 = 32'd9
; 
32'd7017: dataIn1 = 32'd10
; 
32'd7018: dataIn1 = 32'd13
; 
32'd7019: dataIn1 = 32'd15
; 
32'd7020: dataIn1 = 32'd16
; 
32'd7021: dataIn1 = 32'd18
; 
32'd7022: dataIn1 = 32'd19
; 
32'd7023: dataIn1 = 32'd20
; 
32'd7024: dataIn1 = 32'd22
; 
32'd7025: dataIn1 = 32'd23
; 
32'd7026: dataIn1 = 32'd25
; 
32'd7027: dataIn1 = 32'd26
; 
32'd7028: dataIn1 = 32'd28
; 
32'd7029: dataIn1 = 32'd29
; 
32'd7030: dataIn1 = 32'd30
; 
32'd7031: dataIn1 = 32'd0
; 
32'd7032: dataIn1 = 32'd1
; 
32'd7033: dataIn1 = 32'd4
; 
32'd7034: dataIn1 = 32'd5
; 
32'd7035: dataIn1 = 32'd10
; 
32'd7036: dataIn1 = 32'd11
; 
32'd7037: dataIn1 = 32'd12
; 
32'd7038: dataIn1 = 32'd23
; 
32'd7039: dataIn1 = 32'd25
; 
32'd7040: dataIn1 = 32'd27
; 
32'd7041: dataIn1 = 32'd29
; 
32'd7042: dataIn1 = 32'd30
; 
32'd7043: dataIn1 = 32'd31
; 
32'd7044: dataIn1 = 32'd0
; 
32'd7045: dataIn1 = 32'd4
; 
32'd7046: dataIn1 = 32'd7
; 
32'd7047: dataIn1 = 32'd8
; 
32'd7048: dataIn1 = 32'd9
; 
32'd7049: dataIn1 = 32'd12
; 
32'd7050: dataIn1 = 32'd15
; 
32'd7051: dataIn1 = 32'd16
; 
32'd7052: dataIn1 = 32'd18
; 
32'd7053: dataIn1 = 32'd19
; 
32'd7054: dataIn1 = 32'd20
; 
32'd7055: dataIn1 = 32'd22
; 
32'd7056: dataIn1 = 32'd24
; 
32'd7057: dataIn1 = 32'd25
; 
32'd7058: dataIn1 = 32'd26
; 
32'd7059: dataIn1 = 32'd30
; 
32'd7060: dataIn1 = 32'd31
; 
32'd7061: dataIn1 = 32'd0
; 
32'd7062: dataIn1 = 32'd2
; 
32'd7063: dataIn1 = 32'd3
; 
32'd7064: dataIn1 = 32'd5
; 
32'd7065: dataIn1 = 32'd7
; 
32'd7066: dataIn1 = 32'd10
; 
32'd7067: dataIn1 = 32'd13
; 
32'd7068: dataIn1 = 32'd15
; 
32'd7069: dataIn1 = 32'd16
; 
32'd7070: dataIn1 = 32'd17
; 
32'd7071: dataIn1 = 32'd24
; 
32'd7072: dataIn1 = 32'd26
; 
32'd7073: dataIn1 = 32'd27
; 
32'd7074: dataIn1 = 32'd28
; 
32'd7075: dataIn1 = 32'd30
; 
32'd7076: dataIn1 = 32'd2
; 
32'd7077: dataIn1 = 32'd5
; 
32'd7078: dataIn1 = 32'd8
; 
32'd7079: dataIn1 = 32'd10
; 
32'd7080: dataIn1 = 32'd13
; 
32'd7081: dataIn1 = 32'd15
; 
32'd7082: dataIn1 = 32'd16
; 
32'd7083: dataIn1 = 32'd18
; 
32'd7084: dataIn1 = 32'd19
; 
32'd7085: dataIn1 = 32'd20
; 
32'd7086: dataIn1 = 32'd23
; 
32'd7087: dataIn1 = 32'd24
; 
32'd7088: dataIn1 = 32'd29
; 
32'd7089: dataIn1 = 32'd30
; 
32'd7090: dataIn1 = 32'd0
; 
32'd7091: dataIn1 = 32'd2
; 
32'd7092: dataIn1 = 32'd3
; 
32'd7093: dataIn1 = 32'd5
; 
32'd7094: dataIn1 = 32'd7
; 
32'd7095: dataIn1 = 32'd8
; 
32'd7096: dataIn1 = 32'd9
; 
32'd7097: dataIn1 = 32'd12
; 
32'd7098: dataIn1 = 32'd14
; 
32'd7099: dataIn1 = 32'd15
; 
32'd7100: dataIn1 = 32'd17
; 
32'd7101: dataIn1 = 32'd21
; 
32'd7102: dataIn1 = 32'd25
; 
32'd7103: dataIn1 = 32'd26
; 
32'd7104: dataIn1 = 32'd29
; 
32'd7105: dataIn1 = 32'd0
; 
32'd7106: dataIn1 = 32'd5
; 
32'd7107: dataIn1 = 32'd7
; 
32'd7108: dataIn1 = 32'd8
; 
32'd7109: dataIn1 = 32'd9
; 
32'd7110: dataIn1 = 32'd10
; 
32'd7111: dataIn1 = 32'd11
; 
32'd7112: dataIn1 = 32'd14
; 
32'd7113: dataIn1 = 32'd15
; 
32'd7114: dataIn1 = 32'd16
; 
32'd7115: dataIn1 = 32'd17
; 
32'd7116: dataIn1 = 32'd18
; 
32'd7117: dataIn1 = 32'd19
; 
32'd7118: dataIn1 = 32'd20
; 
32'd7119: dataIn1 = 32'd21
; 
32'd7120: dataIn1 = 32'd22
; 
32'd7121: dataIn1 = 32'd24
; 
32'd7122: dataIn1 = 32'd25
; 
32'd7123: dataIn1 = 32'd26
; 
32'd7124: dataIn1 = 32'd28
; 
32'd7125: dataIn1 = 32'd30
; 
32'd7126: dataIn1 = 32'd31
; 
32'd7127: dataIn1 = 32'd0
; 
32'd7128: dataIn1 = 32'd1
; 
32'd7129: dataIn1 = 32'd3
; 
32'd7130: dataIn1 = 32'd5
; 
32'd7131: dataIn1 = 32'd7
; 
32'd7132: dataIn1 = 32'd8
; 
32'd7133: dataIn1 = 32'd9
; 
32'd7134: dataIn1 = 32'd10
; 
32'd7135: dataIn1 = 32'd12
; 
32'd7136: dataIn1 = 32'd13
; 
32'd7137: dataIn1 = 32'd14
; 
32'd7138: dataIn1 = 32'd15
; 
32'd7139: dataIn1 = 32'd17
; 
32'd7140: dataIn1 = 32'd18
; 
32'd7141: dataIn1 = 32'd22
; 
32'd7142: dataIn1 = 32'd23
; 
32'd7143: dataIn1 = 32'd24
; 
32'd7144: dataIn1 = 32'd27
; 
32'd7145: dataIn1 = 32'd28
; 
32'd7146: dataIn1 = 32'd29
; 
32'd7147: dataIn1 = 32'd30
; 
32'd7148: dataIn1 = 32'd31
; 
32'd7149: dataIn1 = 32'd1
; 
32'd7150: dataIn1 = 32'd6
; 
32'd7151: dataIn1 = 32'd7
; 
32'd7152: dataIn1 = 32'd10
; 
32'd7153: dataIn1 = 32'd11
; 
32'd7154: dataIn1 = 32'd14
; 
32'd7155: dataIn1 = 32'd16
; 
32'd7156: dataIn1 = 32'd18
; 
32'd7157: dataIn1 = 32'd25
; 
32'd7158: dataIn1 = 32'd26
; 
32'd7159: dataIn1 = 32'd30
; 
32'd7160: dataIn1 = 32'd0
; 
32'd7161: dataIn1 = 32'd3
; 
32'd7162: dataIn1 = 32'd8
; 
32'd7163: dataIn1 = 32'd10
; 
32'd7164: dataIn1 = 32'd11
; 
32'd7165: dataIn1 = 32'd14
; 
32'd7166: dataIn1 = 32'd16
; 
32'd7167: dataIn1 = 32'd21
; 
32'd7168: dataIn1 = 32'd23
; 
32'd7169: dataIn1 = 32'd26
; 
32'd7170: dataIn1 = 32'd28
; 
32'd7171: dataIn1 = 32'd29
; 
32'd7172: dataIn1 = 32'd31
; 
32'd7173: dataIn1 = 32'd0
; 
32'd7174: dataIn1 = 32'd1
; 
32'd7175: dataIn1 = 32'd3
; 
32'd7176: dataIn1 = 32'd9
; 
32'd7177: dataIn1 = 32'd10
; 
32'd7178: dataIn1 = 32'd12
; 
32'd7179: dataIn1 = 32'd14
; 
32'd7180: dataIn1 = 32'd16
; 
32'd7181: dataIn1 = 32'd23
; 
32'd7182: dataIn1 = 32'd24
; 
32'd7183: dataIn1 = 32'd25
; 
32'd7184: dataIn1 = 32'd27
; 
32'd7185: dataIn1 = 32'd31
; 
32'd7186: dataIn1 = 32'd2
; 
32'd7187: dataIn1 = 32'd5
; 
32'd7188: dataIn1 = 32'd9
; 
32'd7189: dataIn1 = 32'd10
; 
32'd7190: dataIn1 = 32'd11
; 
32'd7191: dataIn1 = 32'd15
; 
32'd7192: dataIn1 = 32'd19
; 
32'd7193: dataIn1 = 32'd26
; 
32'd7194: dataIn1 = 32'd28
; 
32'd7195: dataIn1 = 32'd29
; 
32'd7196: dataIn1 = 32'd30
; 
32'd7197: dataIn1 = 32'd31
; 
32'd7198: dataIn1 = 32'd0
; 
32'd7199: dataIn1 = 32'd1
; 
32'd7200: dataIn1 = 32'd2
; 
32'd7201: dataIn1 = 32'd4
; 
32'd7202: dataIn1 = 32'd5
; 
32'd7203: dataIn1 = 32'd7
; 
32'd7204: dataIn1 = 32'd10
; 
32'd7205: dataIn1 = 32'd11
; 
32'd7206: dataIn1 = 32'd13
; 
32'd7207: dataIn1 = 32'd17
; 
32'd7208: dataIn1 = 32'd20
; 
32'd7209: dataIn1 = 32'd22
; 
32'd7210: dataIn1 = 32'd23
; 
32'd7211: dataIn1 = 32'd28
; 
32'd7212: dataIn1 = 32'd29
; 
32'd7213: dataIn1 = 32'd0
; 
32'd7214: dataIn1 = 32'd3
; 
32'd7215: dataIn1 = 32'd4
; 
32'd7216: dataIn1 = 32'd13
; 
32'd7217: dataIn1 = 32'd14
; 
32'd7218: dataIn1 = 32'd16
; 
32'd7219: dataIn1 = 32'd17
; 
32'd7220: dataIn1 = 32'd21
; 
32'd7221: dataIn1 = 32'd22
; 
32'd7222: dataIn1 = 32'd24
; 
32'd7223: dataIn1 = 32'd28
; 
32'd7224: dataIn1 = 32'd31
; 
32'd7225: dataIn1 = 32'd2
; 
32'd7226: dataIn1 = 32'd3
; 
32'd7227: dataIn1 = 32'd5
; 
32'd7228: dataIn1 = 32'd7
; 
32'd7229: dataIn1 = 32'd8
; 
32'd7230: dataIn1 = 32'd9
; 
32'd7231: dataIn1 = 32'd13
; 
32'd7232: dataIn1 = 32'd15
; 
32'd7233: dataIn1 = 32'd17
; 
32'd7234: dataIn1 = 32'd23
; 
32'd7235: dataIn1 = 32'd26
; 
32'd7236: dataIn1 = 32'd27
; 
32'd7237: dataIn1 = 32'd29
; 
32'd7238: dataIn1 = 32'd30
; 
32'd7239: dataIn1 = 32'd0
; 
32'd7240: dataIn1 = 32'd1
; 
32'd7241: dataIn1 = 32'd3
; 
32'd7242: dataIn1 = 32'd5
; 
32'd7243: dataIn1 = 32'd6
; 
32'd7244: dataIn1 = 32'd7
; 
32'd7245: dataIn1 = 32'd10
; 
32'd7246: dataIn1 = 32'd11
; 
32'd7247: dataIn1 = 32'd12
; 
32'd7248: dataIn1 = 32'd15
; 
32'd7249: dataIn1 = 32'd17
; 
32'd7250: dataIn1 = 32'd18
; 
32'd7251: dataIn1 = 32'd19
; 
32'd7252: dataIn1 = 32'd21
; 
32'd7253: dataIn1 = 32'd24
; 
32'd7254: dataIn1 = 32'd26
; 
32'd7255: dataIn1 = 32'd28
; 
32'd7256: dataIn1 = 32'd29
; 
32'd7257: dataIn1 = 32'd31
; 
32'd7258: dataIn1 = 32'd0
; 
32'd7259: dataIn1 = 32'd2
; 
32'd7260: dataIn1 = 32'd3
; 
32'd7261: dataIn1 = 32'd4
; 
32'd7262: dataIn1 = 32'd12
; 
32'd7263: dataIn1 = 32'd13
; 
32'd7264: dataIn1 = 32'd16
; 
32'd7265: dataIn1 = 32'd17
; 
32'd7266: dataIn1 = 32'd18
; 
32'd7267: dataIn1 = 32'd20
; 
32'd7268: dataIn1 = 32'd22
; 
32'd7269: dataIn1 = 32'd26
; 
32'd7270: dataIn1 = 32'd27
; 
32'd7271: dataIn1 = 32'd31
; 
32'd7272: dataIn1 = 32'd2
; 
32'd7273: dataIn1 = 32'd3
; 
32'd7274: dataIn1 = 32'd5
; 
32'd7275: dataIn1 = 32'd7
; 
32'd7276: dataIn1 = 32'd8
; 
32'd7277: dataIn1 = 32'd9
; 
32'd7278: dataIn1 = 32'd10
; 
32'd7279: dataIn1 = 32'd11
; 
32'd7280: dataIn1 = 32'd12
; 
32'd7281: dataIn1 = 32'd13
; 
32'd7282: dataIn1 = 32'd14
; 
32'd7283: dataIn1 = 32'd16
; 
32'd7284: dataIn1 = 32'd19
; 
32'd7285: dataIn1 = 32'd21
; 
32'd7286: dataIn1 = 32'd22
; 
32'd7287: dataIn1 = 32'd29
; 
32'd7288: dataIn1 = 32'd30
; 
32'd7289: dataIn1 = 32'd31
; 
32'd7290: dataIn1 = 32'd1
; 
32'd7291: dataIn1 = 32'd2
; 
32'd7292: dataIn1 = 32'd5
; 
32'd7293: dataIn1 = 32'd7
; 
32'd7294: dataIn1 = 32'd9
; 
32'd7295: dataIn1 = 32'd10
; 
32'd7296: dataIn1 = 32'd14
; 
32'd7297: dataIn1 = 32'd15
; 
32'd7298: dataIn1 = 32'd16
; 
32'd7299: dataIn1 = 32'd19
; 
32'd7300: dataIn1 = 32'd20
; 
32'd7301: dataIn1 = 32'd21
; 
32'd7302: dataIn1 = 32'd22
; 
32'd7303: dataIn1 = 32'd28
; 
32'd7304: dataIn1 = 32'd31
; 
32'd7305: dataIn1 = 32'd1
; 
32'd7306: dataIn1 = 32'd4
; 
32'd7307: dataIn1 = 32'd5
; 
32'd7308: dataIn1 = 32'd6
; 
32'd7309: dataIn1 = 32'd9
; 
32'd7310: dataIn1 = 32'd10
; 
32'd7311: dataIn1 = 32'd11
; 
32'd7312: dataIn1 = 32'd12
; 
32'd7313: dataIn1 = 32'd13
; 
32'd7314: dataIn1 = 32'd16
; 
32'd7315: dataIn1 = 32'd17
; 
32'd7316: dataIn1 = 32'd18
; 
32'd7317: dataIn1 = 32'd19
; 
32'd7318: dataIn1 = 32'd21
; 
32'd7319: dataIn1 = 32'd22
; 
32'd7320: dataIn1 = 32'd23
; 
32'd7321: dataIn1 = 32'd25
; 
32'd7322: dataIn1 = 32'd26
; 
32'd7323: dataIn1 = 32'd27
; 
32'd7324: dataIn1 = 32'd29
; 
32'd7325: dataIn1 = 32'd30
; 
32'd7326: dataIn1 = 32'd4
; 
32'd7327: dataIn1 = 32'd6
; 
32'd7328: dataIn1 = 32'd8
; 
32'd7329: dataIn1 = 32'd9
; 
32'd7330: dataIn1 = 32'd11
; 
32'd7331: dataIn1 = 32'd16
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd34; 
32'd3: dataIn2 = 32'd83; 
32'd4: dataIn2 = 32'd61; 
32'd5: dataIn2 = 32'd5; 
32'd6: dataIn2 = 32'd34; 
32'd7: dataIn2 = 32'd77; 
32'd8: dataIn2 = 32'd26; 
32'd9: dataIn2 = 32'd99; 
32'd10: dataIn2 = 32'd68; 
32'd11: dataIn2 = 32'd8; 
32'd12: dataIn2 = 32'd49; 
32'd13: dataIn2 = 32'd22; 
32'd14: dataIn2 = 32'd28; 
32'd15: dataIn2 = 32'd62; 
32'd16: dataIn2 = 32'd53; 
32'd17: dataIn2 = 32'd16; 
32'd18: dataIn2 = 32'd53; 
32'd19: dataIn2 = 32'd3; 
32'd20: dataIn2 = 32'd33; 
32'd21: dataIn2 = 32'd35; 
32'd22: dataIn2 = 32'd27; 
32'd23: dataIn2 = 32'd13; 
32'd24: dataIn2 = 32'd56; 
32'd25: dataIn2 = 32'd70; 
32'd26: dataIn2 = 32'd44; 
32'd27: dataIn2 = 32'd12; 
32'd28: dataIn2 = 32'd87; 
32'd29: dataIn2 = 32'd78; 
32'd30: dataIn2 = 32'd29; 
32'd31: dataIn2 = 32'd12; 
32'd32: dataIn2 = 32'd97; 
32'd33: dataIn2 = 32'd48; 
default: 
	dataIn2 = 32'd99999; 
endcase 
32'd170: dataIn2 = 32'd55; 
32'd171: dataIn2 = 32'd74; 
32'd172: dataIn2 = 32'd12; 
32'd173: dataIn2 = 32'd54; 
32'd174: dataIn2 = 32'd35; 
32'd175: dataIn2 = 32'd39; 
32'd176: dataIn2 = 32'd53; 
32'd177: dataIn2 = 32'd16; 
32'd178: dataIn2 = 32'd44; 
32'd179: dataIn2 = 32'd27; 
32'd180: dataIn2 = 32'd96; 
32'd181: dataIn2 = 32'd50; 
32'd182: dataIn2 = 32'd51; 
32'd183: dataIn2 = 32'd29; 
32'd184: dataIn2 = 32'd44; 
32'd185: dataIn2 = 32'd25; 
32'd186: dataIn2 = 32'd23; 
32'd187: dataIn2 = 32'd33; 
32'd188: dataIn2 = 32'd20; 
32'd189: dataIn2 = 32'd77; 
32'd190: dataIn2 = 32'd80; 
32'd191: dataIn2 = 32'd62; 
32'd192: dataIn2 = 32'd19; 
32'd193: dataIn2 = 32'd51; 
32'd194: dataIn2 = 32'd26; 
32'd195: dataIn2 = 32'd91; 
32'd196: dataIn2 = 32'd90; 
32'd197: dataIn2 = 32'd76; 
32'd198: dataIn2 = 32'd85; 
32'd199: dataIn2 = 32'd77; 
32'd200: dataIn2 = 32'd7; 
32'd201: dataIn2 = 32'd21; 
32'd202: dataIn2 = 32'd27; 
32'd203: dataIn2 = 32'd36; 
32'd204: dataIn2 = 32'd74; 
32'd205: dataIn2 = 32'd71; 
32'd206: dataIn2 = 32'd17; 
32'd207: dataIn2 = 32'd90; 
32'd208: dataIn2 = 32'd55; 
32'd209: dataIn2 = 32'd34; 
32'd210: dataIn2 = 32'd55; 
32'd211: dataIn2 = 32'd14; 
32'd212: dataIn2 = 32'd9; 
32'd213: dataIn2 = 32'd76; 
32'd214: dataIn2 = 32'd29; 
32'd215: dataIn2 = 32'd69; 
32'd216: dataIn2 = 32'd29; 
32'd217: dataIn2 = 32'd50; 
32'd218: dataIn2 = 32'd22; 
32'd219: dataIn2 = 32'd87; 
32'd220: dataIn2 = 32'd15; 
32'd221: dataIn2 = 32'd77; 
32'd222: dataIn2 = 32'd20; 
32'd223: dataIn2 = 32'd14; 
32'd224: dataIn2 = 32'd80; 
32'd225: dataIn2 = 32'd35; 
32'd226: dataIn2 = 32'd24; 
32'd227: dataIn2 = 32'd94; 
32'd228: dataIn2 = 32'd68; 
32'd229: dataIn2 = 32'd47; 
32'd230: dataIn2 = 32'd18; 
32'd231: dataIn2 = 32'd95; 
32'd232: dataIn2 = 32'd80; 
32'd233: dataIn2 = 32'd14; 
32'd234: dataIn2 = 32'd9; 
32'd235: dataIn2 = 32'd9; 
32'd236: dataIn2 = 32'd89; 
32'd237: dataIn2 = 32'd84; 
32'd238: dataIn2 = 32'd80; 
32'd239: dataIn2 = 32'd21; 
32'd240: dataIn2 = 32'd43; 
32'd241: dataIn2 = 32'd40; 
32'd242: dataIn2 = 32'd18; 
32'd243: dataIn2 = 32'd60; 
32'd244: dataIn2 = 32'd63; 
32'd245: dataIn2 = 32'd60; 
32'd246: dataIn2 = 32'd14; 
32'd247: dataIn2 = 32'd73; 
32'd248: dataIn2 = 32'd64; 
32'd249: dataIn2 = 32'd56; 
32'd250: dataIn2 = 32'd76; 
32'd251: dataIn2 = 32'd74; 
32'd252: dataIn2 = 32'd15; 
32'd253: dataIn2 = 32'd45; 
32'd254: dataIn2 = 32'd82; 
32'd255: dataIn2 = 32'd5; 
32'd256: dataIn2 = 32'd98; 
32'd257: dataIn2 = 32'd70; 
32'd258: dataIn2 = 32'd72; 
32'd259: dataIn2 = 32'd44; 
32'd260: dataIn2 = 32'd64; 
32'd261: dataIn2 = 32'd84; 
32'd262: dataIn2 = 32'd2; 
32'd263: dataIn2 = 32'd67; 
32'd264: dataIn2 = 32'd8; 
32'd265: dataIn2 = 32'd89; 
32'd266: dataIn2 = 32'd6; 
32'd267: dataIn2 = 32'd78; 
32'd268: dataIn2 = 32'd66; 
32'd269: dataIn2 = 32'd100; 
32'd270: dataIn2 = 32'd73; 
32'd271: dataIn2 = 32'd34; 
32'd272: dataIn2 = 32'd74; 
32'd273: dataIn2 = 32'd1; 
32'd274: dataIn2 = 32'd37; 
32'd275: dataIn2 = 32'd82; 
32'd276: dataIn2 = 32'd19; 
32'd277: dataIn2 = 32'd86; 
32'd278: dataIn2 = 32'd64; 
32'd279: dataIn2 = 32'd11; 
32'd280: dataIn2 = 32'd60; 
32'd281: dataIn2 = 32'd75; 
32'd282: dataIn2 = 32'd39; 
32'd283: dataIn2 = 32'd13; 
32'd284: dataIn2 = 32'd60; 
32'd285: dataIn2 = 32'd52; 
32'd286: dataIn2 = 32'd60; 
32'd287: dataIn2 = 32'd28; 
32'd288: dataIn2 = 32'd17; 
32'd289: dataIn2 = 32'd16; 
32'd290: dataIn2 = 32'd82; 
32'd291: dataIn2 = 32'd46; 
32'd292: dataIn2 = 32'd58; 
32'd293: dataIn2 = 32'd26; 
32'd294: dataIn2 = 32'd6; 
32'd295: dataIn2 = 32'd37; 
32'd296: dataIn2 = 32'd27; 
32'd297: dataIn2 = 32'd8; 
32'd298: dataIn2 = 32'd76; 
32'd299: dataIn2 = 32'd33; 
32'd300: dataIn2 = 32'd63; 
32'd301: dataIn2 = 32'd84; 
32'd302: dataIn2 = 32'd20; 
32'd303: dataIn2 = 32'd75; 
32'd304: dataIn2 = 32'd63; 
32'd305: dataIn2 = 32'd14; 
32'd306: dataIn2 = 32'd35; 
32'd307: dataIn2 = 32'd36; 
32'd308: dataIn2 = 32'd28; 
32'd309: dataIn2 = 32'd40; 
32'd310: dataIn2 = 32'd36; 
32'd311: dataIn2 = 32'd61; 
32'd312: dataIn2 = 32'd78; 
32'd313: dataIn2 = 32'd34; 
32'd314: dataIn2 = 32'd80; 
32'd315: dataIn2 = 32'd45; 
32'd316: dataIn2 = 32'd50; 
32'd317: dataIn2 = 32'd80; 
32'd318: dataIn2 = 32'd41; 
32'd319: dataIn2 = 32'd50; 
32'd320: dataIn2 = 32'd100; 
32'd321: dataIn2 = 32'd98; 
32'd322: dataIn2 = 32'd13; 
32'd323: dataIn2 = 32'd32; 
32'd324: dataIn2 = 32'd51; 
32'd325: dataIn2 = 32'd66; 
32'd326: dataIn2 = 32'd90; 
32'd327: dataIn2 = 32'd61; 
32'd328: dataIn2 = 32'd87; 
32'd329: dataIn2 = 32'd27; 
32'd330: dataIn2 = 32'd88; 
32'd331: dataIn2 = 32'd86; 
32'd332: dataIn2 = 32'd63; 
32'd333: dataIn2 = 32'd6; 
32'd334: dataIn2 = 32'd9; 
32'd335: dataIn2 = 32'd48; 
32'd336: dataIn2 = 32'd64; 
32'd337: dataIn2 = 32'd2; 
32'd338: dataIn2 = 32'd81; 
32'd339: dataIn2 = 32'd2; 
32'd340: dataIn2 = 32'd69; 
32'd341: dataIn2 = 32'd11; 
32'd342: dataIn2 = 32'd79; 
32'd343: dataIn2 = 32'd56; 
32'd344: dataIn2 = 32'd45; 
32'd345: dataIn2 = 32'd29; 
32'd346: dataIn2 = 32'd53; 
32'd347: dataIn2 = 32'd22; 
32'd348: dataIn2 = 32'd6; 
32'd349: dataIn2 = 32'd87; 
32'd350: dataIn2 = 32'd16; 
32'd351: dataIn2 = 32'd55; 
32'd352: dataIn2 = 32'd35; 
32'd353: dataIn2 = 32'd31; 
32'd354: dataIn2 = 32'd92; 
32'd355: dataIn2 = 32'd7; 
32'd356: dataIn2 = 32'd62; 
32'd357: dataIn2 = 32'd81; 
32'd358: dataIn2 = 32'd53; 
32'd359: dataIn2 = 32'd96; 
32'd360: dataIn2 = 32'd100; 
32'd361: dataIn2 = 32'd6; 
32'd362: dataIn2 = 32'd49; 
32'd363: dataIn2 = 32'd84; 
32'd364: dataIn2 = 32'd92; 
32'd365: dataIn2 = 32'd51; 
32'd366: dataIn2 = 32'd13; 
32'd367: dataIn2 = 32'd62; 
32'd368: dataIn2 = 32'd11; 
32'd369: dataIn2 = 32'd96; 
32'd370: dataIn2 = 32'd67; 
32'd371: dataIn2 = 32'd41; 
32'd372: dataIn2 = 32'd37; 
32'd373: dataIn2 = 32'd17; 
32'd374: dataIn2 = 32'd93; 
32'd375: dataIn2 = 32'd50; 
32'd376: dataIn2 = 32'd50; 
32'd377: dataIn2 = 32'd97; 
32'd378: dataIn2 = 32'd25; 
32'd379: dataIn2 = 32'd52; 
32'd380: dataIn2 = 32'd76; 
32'd381: dataIn2 = 32'd61; 
32'd382: dataIn2 = 32'd1; 
32'd383: dataIn2 = 32'd64; 
32'd384: dataIn2 = 32'd88; 
32'd385: dataIn2 = 32'd65; 
32'd386: dataIn2 = 32'd7; 
32'd387: dataIn2 = 32'd68; 
32'd388: dataIn2 = 32'd64; 
32'd389: dataIn2 = 32'd20; 
32'd390: dataIn2 = 32'd99; 
32'd391: dataIn2 = 32'd77; 
32'd392: dataIn2 = 32'd35; 
32'd393: dataIn2 = 32'd46; 
32'd394: dataIn2 = 32'd76; 
32'd395: dataIn2 = 32'd40; 
32'd396: dataIn2 = 32'd26; 
32'd397: dataIn2 = 32'd22; 
32'd398: dataIn2 = 32'd77; 
32'd399: dataIn2 = 32'd8; 
32'd400: dataIn2 = 32'd26; 
32'd401: dataIn2 = 32'd54; 
32'd402: dataIn2 = 32'd75; 
32'd403: dataIn2 = 32'd25; 
32'd404: dataIn2 = 32'd37; 
32'd405: dataIn2 = 32'd96; 
32'd406: dataIn2 = 32'd90; 
32'd407: dataIn2 = 32'd65; 
32'd408: dataIn2 = 32'd24; 
32'd409: dataIn2 = 32'd24; 
32'd410: dataIn2 = 32'd28; 
32'd411: dataIn2 = 32'd98; 
32'd412: dataIn2 = 32'd19; 
32'd413: dataIn2 = 32'd54; 
32'd414: dataIn2 = 32'd16; 
32'd415: dataIn2 = 32'd91; 
32'd416: dataIn2 = 32'd10; 
32'd417: dataIn2 = 32'd8; 
32'd418: dataIn2 = 32'd12; 
32'd419: dataIn2 = 32'd6; 
32'd420: dataIn2 = 32'd34; 
32'd421: dataIn2 = 32'd97; 
32'd422: dataIn2 = 32'd25; 
32'd423: dataIn2 = 32'd44; 
32'd424: dataIn2 = 32'd75; 
32'd425: dataIn2 = 32'd13; 
32'd426: dataIn2 = 32'd66; 
32'd427: dataIn2 = 32'd30; 
32'd428: dataIn2 = 32'd14; 
32'd429: dataIn2 = 32'd94; 
32'd430: dataIn2 = 32'd48; 
32'd431: dataIn2 = 32'd42; 
32'd432: dataIn2 = 32'd95; 
32'd433: dataIn2 = 32'd82; 
32'd434: dataIn2 = 32'd15; 
32'd435: dataIn2 = 32'd6; 
32'd436: dataIn2 = 32'd76; 
32'd437: dataIn2 = 32'd60; 
32'd438: dataIn2 = 32'd20; 
32'd439: dataIn2 = 32'd0; 
32'd440: dataIn2 = 32'd48; 
32'd441: dataIn2 = 32'd93; 
32'd442: dataIn2 = 32'd99; 
32'd443: dataIn2 = 32'd89; 
32'd444: dataIn2 = 32'd72; 
32'd445: dataIn2 = 32'd29; 
32'd446: dataIn2 = 32'd4; 
32'd447: dataIn2 = 32'd86; 
32'd448: dataIn2 = 32'd78; 
32'd449: dataIn2 = 32'd14; 
32'd450: dataIn2 = 32'd9; 
32'd451: dataIn2 = 32'd50; 
32'd452: dataIn2 = 32'd25; 
32'd453: dataIn2 = 32'd70; 
32'd454: dataIn2 = 32'd51; 
32'd455: dataIn2 = 32'd44; 
32'd456: dataIn2 = 32'd77; 
32'd457: dataIn2 = 32'd32; 
32'd458: dataIn2 = 32'd93; 
32'd459: dataIn2 = 32'd95; 
32'd460: dataIn2 = 32'd75; 
32'd461: dataIn2 = 32'd20; 
32'd462: dataIn2 = 32'd4; 
32'd463: dataIn2 = 32'd62; 
32'd464: dataIn2 = 32'd2; 
32'd465: dataIn2 = 32'd33; 
32'd466: dataIn2 = 32'd23; 
32'd467: dataIn2 = 32'd11; 
32'd468: dataIn2 = 32'd75; 
32'd469: dataIn2 = 32'd47; 
32'd470: dataIn2 = 32'd87; 
32'd471: dataIn2 = 32'd63; 
32'd472: dataIn2 = 32'd89; 
32'd473: dataIn2 = 32'd41; 
32'd474: dataIn2 = 32'd3; 
32'd475: dataIn2 = 32'd31; 
32'd476: dataIn2 = 32'd15; 
32'd477: dataIn2 = 32'd71; 
32'd478: dataIn2 = 32'd45; 
32'd479: dataIn2 = 32'd46; 
32'd480: dataIn2 = 32'd7; 
32'd481: dataIn2 = 32'd62; 
32'd482: dataIn2 = 32'd81; 
32'd483: dataIn2 = 32'd38; 
32'd484: dataIn2 = 32'd80; 
32'd485: dataIn2 = 32'd51; 
32'd486: dataIn2 = 32'd35; 
32'd487: dataIn2 = 32'd81; 
32'd488: dataIn2 = 32'd90; 
32'd489: dataIn2 = 32'd99; 
32'd490: dataIn2 = 32'd51; 
32'd491: dataIn2 = 32'd16; 
32'd492: dataIn2 = 32'd29; 
32'd493: dataIn2 = 32'd79; 
32'd494: dataIn2 = 32'd52; 
32'd495: dataIn2 = 32'd93; 
32'd496: dataIn2 = 32'd39; 
32'd497: dataIn2 = 32'd91; 
32'd498: dataIn2 = 32'd13; 
32'd499: dataIn2 = 32'd74; 
32'd500: dataIn2 = 32'd3; 
32'd501: dataIn2 = 32'd71; 
32'd502: dataIn2 = 32'd75; 
32'd503: dataIn2 = 32'd44; 
32'd504: dataIn2 = 32'd61; 
32'd505: dataIn2 = 32'd52; 
32'd506: dataIn2 = 32'd80; 
32'd507: dataIn2 = 32'd0; 
32'd508: dataIn2 = 32'd34; 
32'd509: dataIn2 = 32'd62; 
32'd510: dataIn2 = 32'd33; 
32'd511: dataIn2 = 32'd90; 
32'd512: dataIn2 = 32'd88; 
32'd513: dataIn2 = 32'd52; 
32'd514: dataIn2 = 32'd98; 
32'd515: dataIn2 = 32'd2; 
32'd516: dataIn2 = 32'd45; 
32'd517: dataIn2 = 32'd20; 
32'd518: dataIn2 = 32'd67; 
32'd519: dataIn2 = 32'd44; 
32'd520: dataIn2 = 32'd98; 
32'd521: dataIn2 = 32'd13; 
32'd522: dataIn2 = 32'd63; 
32'd523: dataIn2 = 32'd94; 
32'd524: dataIn2 = 32'd12; 
32'd525: dataIn2 = 32'd100; 
32'd526: dataIn2 = 32'd48; 
32'd527: dataIn2 = 32'd27; 
32'd528: dataIn2 = 32'd24; 
32'd529: dataIn2 = 32'd12; 
32'd530: dataIn2 = 32'd98; 
32'd531: dataIn2 = 32'd86; 
32'd532: dataIn2 = 32'd29; 
32'd533: dataIn2 = 32'd15; 
32'd534: dataIn2 = 32'd37; 
32'd535: dataIn2 = 32'd36; 
32'd536: dataIn2 = 32'd88; 
32'd537: dataIn2 = 32'd74; 
32'd538: dataIn2 = 32'd69; 
32'd539: dataIn2 = 32'd94; 
32'd540: dataIn2 = 32'd35; 
32'd541: dataIn2 = 32'd46; 
32'd542: dataIn2 = 32'd85; 
32'd543: dataIn2 = 32'd28; 
32'd544: dataIn2 = 32'd10; 
32'd545: dataIn2 = 32'd93; 
32'd546: dataIn2 = 32'd41; 
32'd547: dataIn2 = 32'd91; 
32'd548: dataIn2 = 32'd73; 
32'd549: dataIn2 = 32'd27; 
32'd550: dataIn2 = 32'd49; 
32'd551: dataIn2 = 32'd40; 
32'd552: dataIn2 = 32'd97; 
32'd553: dataIn2 = 32'd22; 
32'd554: dataIn2 = 32'd3; 
32'd555: dataIn2 = 32'd76; 
32'd556: dataIn2 = 32'd77; 
32'd557: dataIn2 = 32'd3; 
32'd558: dataIn2 = 32'd81; 
32'd559: dataIn2 = 32'd72; 
32'd560: dataIn2 = 32'd18; 
32'd561: dataIn2 = 32'd64; 
32'd562: dataIn2 = 32'd78; 
32'd563: dataIn2 = 32'd62; 
32'd564: dataIn2 = 32'd97; 
32'd565: dataIn2 = 32'd39; 
32'd566: dataIn2 = 32'd96; 
32'd567: dataIn2 = 32'd66; 
32'd568: dataIn2 = 32'd49; 
32'd569: dataIn2 = 32'd51; 
32'd570: dataIn2 = 32'd80; 
32'd571: dataIn2 = 32'd78; 
32'd572: dataIn2 = 32'd83; 
32'd573: dataIn2 = 32'd93; 
32'd574: dataIn2 = 32'd94; 
32'd575: dataIn2 = 32'd46; 
32'd576: dataIn2 = 32'd35; 
32'd577: dataIn2 = 32'd78; 
32'd578: dataIn2 = 32'd67; 
32'd579: dataIn2 = 32'd1; 
32'd580: dataIn2 = 32'd92; 
32'd581: dataIn2 = 32'd83; 
32'd582: dataIn2 = 32'd32; 
32'd583: dataIn2 = 32'd6; 
32'd584: dataIn2 = 32'd69; 
32'd585: dataIn2 = 32'd35; 
32'd586: dataIn2 = 32'd55; 
32'd587: dataIn2 = 32'd10; 
32'd588: dataIn2 = 32'd9; 
32'd589: dataIn2 = 32'd23; 
32'd590: dataIn2 = 32'd90; 
32'd591: dataIn2 = 32'd63; 
32'd592: dataIn2 = 32'd42; 
32'd593: dataIn2 = 32'd79; 
32'd594: dataIn2 = 32'd34; 
32'd595: dataIn2 = 32'd80; 
32'd596: dataIn2 = 32'd22; 
32'd597: dataIn2 = 32'd50; 
32'd598: dataIn2 = 32'd20; 
32'd599: dataIn2 = 32'd34; 
32'd600: dataIn2 = 32'd81; 
32'd601: dataIn2 = 32'd42; 
32'd602: dataIn2 = 32'd53; 
32'd603: dataIn2 = 32'd50; 
32'd604: dataIn2 = 32'd13; 
32'd605: dataIn2 = 32'd27; 
32'd606: dataIn2 = 32'd21; 
32'd607: dataIn2 = 32'd93; 
32'd608: dataIn2 = 32'd97; 
32'd609: dataIn2 = 32'd82; 
32'd610: dataIn2 = 32'd19; 
32'd611: dataIn2 = 32'd9; 
32'd612: dataIn2 = 32'd35; 
32'd613: dataIn2 = 32'd91; 
32'd614: dataIn2 = 32'd7; 
32'd615: dataIn2 = 32'd1; 
32'd616: dataIn2 = 32'd81; 
32'd617: dataIn2 = 32'd17; 
32'd618: dataIn2 = 32'd34; 
32'd619: dataIn2 = 32'd28; 
32'd620: dataIn2 = 32'd83; 
32'd621: dataIn2 = 32'd8; 
32'd622: dataIn2 = 32'd81; 
32'd623: dataIn2 = 32'd3; 
32'd624: dataIn2 = 32'd0; 
32'd625: dataIn2 = 32'd31; 
32'd626: dataIn2 = 32'd34; 
32'd627: dataIn2 = 32'd40; 
32'd628: dataIn2 = 32'd70; 
32'd629: dataIn2 = 32'd11; 
32'd630: dataIn2 = 32'd14; 
32'd631: dataIn2 = 32'd7; 
32'd632: dataIn2 = 32'd77; 
32'd633: dataIn2 = 32'd52; 
32'd634: dataIn2 = 32'd25; 
32'd635: dataIn2 = 32'd39; 
32'd636: dataIn2 = 32'd58; 
32'd637: dataIn2 = 32'd92; 
32'd638: dataIn2 = 32'd27; 
32'd639: dataIn2 = 32'd27; 
32'd640: dataIn2 = 32'd56; 
32'd641: dataIn2 = 32'd11; 
32'd642: dataIn2 = 32'd19; 
32'd643: dataIn2 = 32'd23; 
32'd644: dataIn2 = 32'd90; 
32'd645: dataIn2 = 32'd46; 
32'd646: dataIn2 = 32'd59; 
32'd647: dataIn2 = 32'd4; 
32'd648: dataIn2 = 32'd50; 
32'd649: dataIn2 = 32'd33; 
32'd650: dataIn2 = 32'd21; 
32'd651: dataIn2 = 32'd76; 
32'd652: dataIn2 = 32'd5; 
32'd653: dataIn2 = 32'd69; 
32'd654: dataIn2 = 32'd27; 
32'd655: dataIn2 = 32'd4; 
32'd656: dataIn2 = 32'd51; 
32'd657: dataIn2 = 32'd1; 
32'd658: dataIn2 = 32'd65; 
32'd659: dataIn2 = 32'd1; 
32'd660: dataIn2 = 32'd98; 
32'd661: dataIn2 = 32'd59; 
32'd662: dataIn2 = 32'd80; 
32'd663: dataIn2 = 32'd62; 
32'd664: dataIn2 = 32'd33; 
32'd665: dataIn2 = 32'd21; 
32'd666: dataIn2 = 32'd90; 
32'd667: dataIn2 = 32'd30; 
32'd668: dataIn2 = 32'd85; 
32'd669: dataIn2 = 32'd85; 
32'd670: dataIn2 = 32'd95; 
32'd671: dataIn2 = 32'd25; 
32'd672: dataIn2 = 32'd35; 
32'd673: dataIn2 = 32'd39; 
32'd674: dataIn2 = 32'd8; 
32'd675: dataIn2 = 32'd98; 
32'd676: dataIn2 = 32'd47; 
32'd677: dataIn2 = 32'd88; 
32'd678: dataIn2 = 32'd12; 
32'd679: dataIn2 = 32'd12; 
32'd680: dataIn2 = 32'd94; 
32'd681: dataIn2 = 32'd50; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("hht2_32_50.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
